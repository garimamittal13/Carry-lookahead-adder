.include TSMC_180nm.txt  

.param SUPPLY=1.8
.param LAMBDA=0.09u
.param width_N={5*LAMBDA}     
.param width_P={2*width_N}     
.global gnd vdd  
Vdd vdd gnd 'SUPPLY'

.subckt inv in out vdd gnd
M1 out in gnd gnd CMOSN W={width_N} L={2*LAMBDA}
+ AS={5*width_N*LAMBDA} PS={10*LAMBDA+2*width_N} AD={5*width_N*LAMBDA} PD={10*LAMBDA+2*width_N}
M2 out in vdd vdd CMOSP W={width_P} L={2*LAMBDA}
+ AS={5*width_P*LAMBDA} PS={10*LAMBDA+2*width_P} AD={5*width_P*LAMBDA} PD={10*LAMBDA+2*width_P}
.ends inv

.subckt and A B Y vdd gnd
M1 out A vdd vdd CMOSP W={width_P} L={2*LAMBDA}
+ AS={5*width_P*LAMBDA} PS={10*LAMBDA+2*width_P} AD={5*width_P*LAMBDA} PD={10*LAMBDA+2*width_P}
M2 out B vdd vdd CMOSP W={width_P} L={2*LAMBDA}
+ AS={5*width_P*LAMBDA} PS={10*LAMBDA+2*width_P} AD={5*width_P*LAMBDA} PD={10*LAMBDA+2*width_P}
M3 out A C C CMOSN W={2*width_N} L={2*LAMBDA}
+ AS={5*2*width_N*LAMBDA} PS={10*LAMBDA+2*2*width_N} AD={5*2*width_N*LAMBDA} PD={10*2*LAMBDA+2*width_N}
M4 C B gnd gnd CMOSN W={2*width_N} L={2*LAMBDA}
+ AS={5*2*width_N*LAMBDA} PS={10*LAMBDA+2*2*width_N} AD={5*2*width_N*LAMBDA} PD={10*LAMBDA+2*2*width_N}
Xinv out Y vdd gnd inv
.ends and

.subckt or A B Y vdd gnd
M1 C A vdd vdd CMOSP W={2*width_P} L={2*LAMBDA}
+ AS={5*2*width_P*LAMBDA} PS={10*LAMBDA+2*2*width_P} AD={5*2*width_P*LAMBDA} PD={10*LAMBDA+2*2*width_P}
M2 out B C C CMOSP W={2*width_P} L={2*LAMBDA}
+ AS={5*2*width_P*LAMBDA} PS={10*LAMBDA+2*2*width_P} AD={5*2*width_P*LAMBDA} PD={10*LAMBDA+2*2*width_P}
M3 out A gnd gnd CMOSN W={width_N} L={2*LAMBDA}
+ AS={5*width_N*LAMBDA} PS={10*LAMBDA+2*width_N} AD={5*width_N*LAMBDA} PD={10*LAMBDA+2*width_N}
M4 out B gnd gnd CMOSN W={width_N} L={2*LAMBDA}
+ AS={5*width_N*LAMBDA} PS={10*LAMBDA+2*width_N} AD={5*width_N*LAMBDA} PD={10*LAMBDA+2*width_N}
Xinv out Y vdd gnd inv
.ends or

*C0, A0, B0, A1, B1, A2, B2, A3, B3 will be given
*have to find S0, S1, S2, S3, Cout

.subckt sum A B Y vdd gnd
Xa A Anot vdd gnd inv
Xb B Bnot vdd gnd inv
X1 A Bnot O1 vdd gnd and
X2 Anot B O2 vdd gnd and
X3 O1 O2 Y vdd gnd or
.ends sum

.subckt generate A B Y vdd gnd
Xg A B Y vdd gnd and
.ends generate

.subckt propagate A B Y vdd gnd
Xp A B Y vdd gnd sum
.ends propagate

Xp0 A0 B0 P0 vdd gnd propagate
Xp1 A1 B1 P1 vdd gnd propagate
Xp2 A2 B2 P2 vdd gnd propagate
Xp3 A3 B3 P3 vdd gnd propagate
Xg0 A0 B0 G0 vdd gnd generate
Xg1 A1 B1 G1 vdd gnd generate
Xg2 A2 B2 G2 vdd gnd generate
Xg3 A3 B3 G3 vdd gnd generate

X1 P0 C0 X0 vdd gnd and
XC1 G0 X0 C1 vdd gnd or

X2 P1 G0 O1 vdd gnd and
X3 P1 X0 O2 vdd gnd and
X4 O1 O2 O3 vdd gnd or
XC2 G1 O3 C2 vdd gnd or

X5 P2 G1 O4 vdd gnd and
X6 O1 P2 O5 vdd gnd and
X7 P2 O2 O6 vdd gnd and
X8 O5 O4 O7 vdd gnd or
X9 O6 O7 O8 vdd gnd or
XC3 G2 O8 C3 vdd gnd or

X10 P3 G2 O9 vdd gnd and
X11 O4 P3 O10 vdd gnd and
X12 O5 P3 O11 vdd gnd and
X13 O6 P3 O12 vdd gnd and
X14 G3 O9 O13 vdd gnd or
X15 O13 O10 O14 vdd gnd or
X16 O14 O11 O15 vdd gnd or

XCout O15 O12 C4 vdd gnd or
Xs0 P0 C0 S0 vdd gnd sum
Xs1 P1 C1 S1 vdd gnd sum
Xs2 P2 C2 S2 vdd gnd sum
Xs3 P3 C3 S3 vdd gnd sum

* Clock and Data Input Signals
Vc C0 gnd dc 0
Va0 A0 gnd dc 0
Va1 A1 gnd dc 1.8
Va2 A2 gnd dc 1.8
Va3 a3 gnd dc 1.8
Vb0 b0 gnd dc 1.8
Vb1 B1 gnd dc 0
Vb2 B2 gnd PULSE(0 'SUPPLY' 0 0.1n 0.1n 10n 20n)
Vb3 b3 gnd dc 0

.tran 1n 35n 15n
.measure tran tpd_rise
+ TRIG v(b2) VAL='SUPPLY/2' RISE=1
+ TARG v(s3) VAL='SUPPLY/2' FALL=1
.measure tran tpd_fall
+ TRIG v(b2) VAL='SUPPLY/2' FALL=1
+ TARG v(s3) VAL='SUPPLY/2' RISE=1
.measure tran total_prop_delay param='(tpd_rise+tpd_fall)/2'

* Control Block for Plotting
.control
run
set color0=white ** color0 is used to set the background of the plot (manual sec:17.7)
set color1=black ** color1 is used to set the grid color of the plot (manual sec:17.7)
set curplottitle= Garima_2023102069
plot V(S0) v(s1)+2 v(s2)+4 v(s3)+6 v(C4)+8
.endc

.end
