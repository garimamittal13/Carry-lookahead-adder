.include TSMC_180nm.txt  

.param SUPPLY=1.8
.param LAMBDA=0.09u
.param width_N={5*LAMBDA}     
.param width_P={10*LAMBDA}     
.global gnd vdd  
Vdd vdd gnd 'SUPPLY'

.subckt inv in out vdd gnd
M1 out in gnd gnd CMOSN W={width_N} L={2*LAMBDA}
+ AS={5*width_N*LAMBDA} PS={10*LAMBDA+2*width_N} AD={5*width_N*LAMBDA} PD={10*LAMBDA+2*width_N}
M2 out in vdd vdd CMOSP W={width_P} L={2*LAMBDA}
+ AS={5*width_P*LAMBDA} PS={10*LAMBDA+2*width_P} AD={5*width_P*LAMBDA} PD={10*LAMBDA+2*width_P}
.ends inv

.subckt and A B Y vdd gnd
M1 out A vdd vdd CMOSP W={width_P} L={2*LAMBDA}
+ AS={5*width_P*LAMBDA} PS={10*LAMBDA+2*width_P} AD={5*width_P*LAMBDA} PD={10*LAMBDA+2*width_P}
M2 out B vdd vdd CMOSP W={width_P} L={2*LAMBDA}
+ AS={5*width_P*LAMBDA} PS={10*LAMBDA+2*width_P} AD={5*width_P*LAMBDA} PD={10*LAMBDA+2*width_P}
M3 out A C C CMOSN W={2*width_N} L={2*LAMBDA}
+ AS={5*2*width_N*LAMBDA} PS={10*LAMBDA+2*2*width_N} AD={5*2*width_N*LAMBDA} PD={10*2*LAMBDA+2*width_N}
M4 C B gnd gnd CMOSN W={2*width_N} L={2*LAMBDA}
+ AS={5*2*width_N*LAMBDA} PS={10*LAMBDA+2*2*width_N} AD={5*2*width_N*LAMBDA} PD={10*LAMBDA+2*2*width_N}
Xinv out Y vdd gnd inv
.ends and

.subckt or A B Y vdd gnd
M1 C A vdd vdd CMOSP W={2*width_P} L={2*LAMBDA}
+ AS={5*2*width_P*LAMBDA} PS={10*LAMBDA+2*2*width_P} AD={5*2*width_P*LAMBDA} PD={10*LAMBDA+2*2*width_P}
M2 out B C C CMOSP W={2*width_P} L={2*LAMBDA}
+ AS={5*2*width_P*LAMBDA} PS={10*LAMBDA+2*2*width_P} AD={5*2*width_P*LAMBDA} PD={10*LAMBDA+2*2*width_P}
M3 out A gnd gnd CMOSN W={width_N} L={2*LAMBDA}
+ AS={5*width_N*LAMBDA} PS={10*LAMBDA+2*width_N} AD={5*width_N*LAMBDA} PD={10*LAMBDA+2*width_N}
M4 out B gnd gnd CMOSN W={width_N} L={2*LAMBDA}
+ AS={5*width_N*LAMBDA} PS={10*LAMBDA+2*width_N} AD={5*width_N*LAMBDA} PD={10*LAMBDA+2*width_N}
Xinv out Y vdd gnd inv
.ends or

*C0, A0, B0, A1, B1, A2, B2, A3, B3 will be given
*have to find S0, S1, S2, S3, Cout
X1 P0 C0 X0 vdd gnd and
XC1 G0 X0 C1 vdd gnd or

X2 P1 G0 O1 vdd gnd and
X3 P1 X0 O2 vdd gnd and
X4 O1 O2 O3 vdd gnd or
XC2 G1 O3 C2 vdd gnd or

X5 P2 G1 O4 vdd gnd and
X6 O1 P2 O5 vdd gnd and
X7 P2 O2 O6 vdd gnd and
X8 O5 O4 O7 vdd gnd or
X9 O6 O7 O8 vdd gnd or
XC3 G2 O8 C3 vdd gnd or

X10 P3 G2 O9 vdd gnd and
X11 O4 P3 O10 vdd gnd and
X12 O5 P3 O11 vdd gnd and
X13 O6 P3 O12 vdd gnd and
X14 G3 O9 O13 vdd gnd or
X15 O13 O10 O14 vdd gnd or
X16 O14 O11 O15 vdd gnd or
XCout O15 O12 C4 vdd gnd or

VX1 p0 gnd 1.8
VX2 p1 gnd pulse 0 1.8 0ns 100ps 100ps 10ns 20ns
VX3 p2 gnd 0
VX4 p3 gnd pulse 0 1.8 0ns 100ps 100ps 15ns 30ns
VX11 g0 gnd pulse 0 1.8 0ns 100ps 100ps 10ns 20ns
VX21 g1 gnd 1.8
VX31 g2 gnd pulse 0 1.8 0ns 100ps 100ps 5ns 10ns
VX41 g3 gnd 0
VX0 c0 gnd 0

.tran 0.1n 30n
.control
run
set color0=white ** color0 is used to set the background of the plot (manual sec:17.7)
set color1=black ** color1 is used to set the grid color of the plot (manual sec:17.7)
set curplottitle= Garima_2023102069
plot V(c1)+2 v(p0)+4 v(g0)+6 
plot V(c2)+2 v(p1)+4 v(g1)+6 
plot V(c3)+2 v(p2)+4 v(g2)+6 
plot V(c4)+2 v(p3)+4 v(g3)+6 
.endc

.end
