magic
tech scmos
timestamp 1732053369
<< nwell >>
rect -3297 -556 -3265 -523
rect -3245 -556 -3221 -523
rect -3857 -597 -3825 -564
rect -3805 -597 -3781 -564
rect -3167 -569 -3133 -543
rect -2298 -547 -2266 -514
rect -2246 -547 -2222 -514
rect -1668 -526 -1636 -493
rect -1616 -526 -1592 -493
rect -2168 -560 -2134 -534
rect -1538 -539 -1504 -513
rect -3727 -610 -3693 -584
rect -3280 -792 -3246 -766
rect -3234 -782 -3200 -757
rect -3186 -785 -3152 -759
rect -2559 -766 -2525 -740
rect -2513 -756 -2479 -731
rect -2465 -759 -2431 -733
rect -1937 -748 -1903 -722
rect -1891 -738 -1857 -713
rect -1843 -741 -1809 -715
rect -3280 -848 -3246 -822
rect -3232 -848 -3198 -823
rect -3184 -851 -3150 -825
rect -3126 -828 -3092 -790
rect -3077 -825 -3043 -799
rect -2559 -822 -2525 -796
rect -2511 -822 -2477 -797
rect -2463 -825 -2429 -799
rect -2405 -802 -2371 -764
rect -2356 -799 -2322 -773
rect -1937 -804 -1903 -778
rect -1889 -804 -1855 -779
rect -1841 -807 -1807 -781
rect -1783 -784 -1749 -746
rect -1734 -781 -1700 -755
rect -3825 -1038 -3791 -1012
rect -3779 -1028 -3745 -1003
rect -3731 -1031 -3697 -1005
rect -3825 -1094 -3791 -1068
rect -3777 -1094 -3743 -1069
rect -3729 -1097 -3695 -1071
rect -3671 -1074 -3637 -1036
rect -3622 -1071 -3588 -1045
rect -2439 -1134 -2405 -1109
rect -2391 -1137 -2357 -1111
rect -2300 -1193 -2266 -1155
rect -2251 -1190 -2217 -1164
rect -2440 -1257 -2406 -1232
rect -2392 -1260 -2358 -1234
rect -2924 -1290 -2890 -1265
rect -2876 -1293 -2842 -1267
rect -4310 -1345 -4278 -1312
rect -4258 -1345 -4234 -1312
rect -4180 -1358 -4146 -1332
rect -2792 -1338 -2758 -1300
rect -2743 -1335 -2709 -1309
rect -2124 -1313 -2090 -1275
rect -2075 -1310 -2041 -1284
rect -1939 -1304 -1905 -1266
rect -1890 -1301 -1856 -1275
rect -1830 -1301 -1798 -1268
rect -1778 -1301 -1754 -1268
rect -1700 -1314 -1666 -1288
rect -3496 -1407 -3462 -1382
rect -3448 -1410 -3414 -1384
rect -2925 -1396 -2891 -1371
rect -2877 -1399 -2843 -1373
rect -2676 -1377 -2642 -1339
rect -2627 -1374 -2593 -1348
rect -2435 -1380 -2401 -1355
rect -2387 -1383 -2353 -1357
rect -3370 -1481 -3336 -1443
rect -3321 -1478 -3287 -1452
rect -3255 -1471 -3221 -1433
rect -2788 -1440 -2754 -1402
rect -2739 -1437 -2705 -1411
rect -2301 -1437 -2267 -1399
rect -2252 -1434 -2218 -1408
rect -3206 -1468 -3172 -1442
rect -3830 -1525 -3796 -1500
rect -3782 -1528 -3748 -1502
rect -3726 -1529 -3692 -1491
rect -3677 -1526 -3643 -1500
rect -3491 -1516 -3457 -1491
rect -2921 -1493 -2887 -1468
rect -3443 -1519 -3409 -1493
rect -2873 -1496 -2839 -1470
rect -2436 -1508 -2402 -1483
rect -2388 -1511 -2354 -1485
rect -4276 -1656 -4244 -1623
rect -4224 -1656 -4200 -1623
rect -3827 -1628 -3793 -1602
rect -3781 -1618 -3747 -1593
rect -3733 -1621 -3699 -1595
rect -3475 -1626 -3441 -1600
rect -3429 -1616 -3395 -1591
rect -3381 -1619 -3347 -1593
rect -4146 -1669 -4112 -1643
rect -3827 -1684 -3793 -1658
rect -3779 -1684 -3745 -1659
rect -3731 -1687 -3697 -1661
rect -3673 -1664 -3639 -1626
rect -3624 -1661 -3590 -1635
rect -3475 -1682 -3441 -1656
rect -3427 -1682 -3393 -1657
rect -3379 -1685 -3345 -1659
rect -3321 -1662 -3287 -1624
rect -2914 -1626 -2880 -1600
rect -2868 -1616 -2834 -1591
rect -2820 -1619 -2786 -1593
rect -2239 -1607 -2205 -1581
rect -2193 -1597 -2159 -1572
rect -2145 -1600 -2111 -1574
rect -3272 -1659 -3238 -1633
rect -2914 -1682 -2880 -1656
rect -2866 -1682 -2832 -1657
rect -2818 -1685 -2784 -1659
rect -2760 -1662 -2726 -1624
rect -2711 -1659 -2677 -1633
rect -2239 -1663 -2205 -1637
rect -2191 -1663 -2157 -1638
rect -2143 -1666 -2109 -1640
rect -2085 -1643 -2051 -1605
rect -2036 -1640 -2002 -1614
rect -2204 -1742 -2170 -1717
rect -2156 -1745 -2122 -1719
rect -3811 -1793 -3777 -1768
rect -3763 -1796 -3729 -1770
rect -3424 -1773 -3390 -1748
rect -3376 -1776 -3342 -1750
rect -2874 -1772 -2840 -1747
rect -2826 -1775 -2792 -1749
rect -4257 -1847 -4225 -1814
rect -4205 -1847 -4181 -1814
rect -4127 -1860 -4093 -1834
rect -2958 -1850 -2926 -1817
rect -2906 -1850 -2882 -1817
rect -2828 -1863 -2794 -1837
rect -2720 -1846 -2688 -1813
rect -2668 -1846 -2644 -1813
rect -2590 -1859 -2556 -1833
rect -2271 -1835 -2239 -1802
rect -2219 -1835 -2195 -1802
rect -2141 -1848 -2107 -1822
rect -1954 -1828 -1922 -1795
rect -1902 -1828 -1878 -1795
rect -1824 -1841 -1790 -1815
rect -3633 -2008 -3601 -1975
rect -3581 -2008 -3557 -1975
rect -3503 -2021 -3469 -1995
rect -3334 -1999 -3302 -1966
rect -3282 -1999 -3258 -1966
rect -3204 -2012 -3170 -1986
<< n_field_implant >>
rect -3211 -556 -3187 -523
rect -2212 -547 -2188 -514
rect -1582 -526 -1558 -493
rect -3771 -597 -3747 -564
rect -1744 -1301 -1720 -1268
rect -4224 -1345 -4200 -1312
rect -4190 -1656 -4166 -1623
rect -4171 -1847 -4147 -1814
rect -2872 -1850 -2848 -1817
rect -2634 -1846 -2610 -1813
rect -2185 -1835 -2161 -1802
rect -1868 -1828 -1844 -1795
rect -3547 -2008 -3523 -1975
rect -3248 -1999 -3224 -1966
<< ntransistor >>
rect -3286 -574 -3284 -569
rect -3846 -615 -3844 -610
rect -3242 -585 -3240 -575
rect -3234 -585 -3232 -575
rect -3200 -585 -3198 -575
rect -3192 -585 -3190 -575
rect -2287 -565 -2285 -560
rect -1657 -544 -1655 -539
rect -2243 -576 -2241 -566
rect -2235 -576 -2233 -566
rect -2201 -576 -2199 -566
rect -2193 -576 -2191 -566
rect -1613 -555 -1611 -545
rect -1605 -555 -1603 -545
rect -1571 -555 -1569 -545
rect -1563 -555 -1561 -545
rect -1526 -553 -1524 -548
rect -2156 -574 -2154 -569
rect -3155 -583 -3153 -578
rect -3802 -626 -3800 -616
rect -3794 -626 -3792 -616
rect -3760 -626 -3758 -616
rect -3752 -626 -3750 -616
rect -3715 -624 -3713 -619
rect -1925 -762 -1923 -757
rect -1880 -761 -1878 -751
rect -1870 -761 -1868 -751
rect -1831 -755 -1829 -750
rect -2547 -780 -2545 -775
rect -2502 -779 -2500 -769
rect -2492 -779 -2490 -769
rect -2453 -773 -2451 -768
rect -3268 -806 -3266 -801
rect -3223 -805 -3221 -795
rect -3213 -805 -3211 -795
rect -3174 -799 -3172 -794
rect -3268 -862 -3266 -857
rect -3065 -839 -3063 -834
rect -2547 -836 -2545 -831
rect -2344 -813 -2342 -808
rect -2394 -821 -2392 -816
rect -2384 -821 -2382 -816
rect -1925 -818 -1923 -813
rect -1722 -795 -1720 -790
rect -1772 -803 -1770 -798
rect -1762 -803 -1760 -798
rect -1878 -827 -1876 -817
rect -1868 -827 -1866 -817
rect -1829 -821 -1827 -816
rect -3115 -847 -3113 -842
rect -3105 -847 -3103 -842
rect -2500 -845 -2498 -835
rect -2490 -845 -2488 -835
rect -2451 -839 -2449 -834
rect -3221 -871 -3219 -861
rect -3211 -871 -3209 -861
rect -3172 -865 -3170 -860
rect -3813 -1052 -3811 -1047
rect -3768 -1051 -3766 -1041
rect -3758 -1051 -3756 -1041
rect -3719 -1045 -3717 -1040
rect -3813 -1108 -3811 -1103
rect -3610 -1085 -3608 -1080
rect -3660 -1093 -3658 -1088
rect -3650 -1093 -3648 -1088
rect -3766 -1117 -3764 -1107
rect -3756 -1117 -3754 -1107
rect -3717 -1111 -3715 -1106
rect -2428 -1157 -2426 -1147
rect -2418 -1157 -2416 -1147
rect -2379 -1151 -2377 -1146
rect -2239 -1204 -2237 -1199
rect -2289 -1212 -2287 -1207
rect -2279 -1212 -2277 -1207
rect -2429 -1280 -2427 -1270
rect -2419 -1280 -2417 -1270
rect -2380 -1274 -2378 -1269
rect -2913 -1313 -2911 -1303
rect -2903 -1313 -2901 -1303
rect -2864 -1307 -2862 -1302
rect -1878 -1315 -1876 -1310
rect -2063 -1324 -2061 -1319
rect -1928 -1323 -1926 -1318
rect -1918 -1323 -1916 -1318
rect -1819 -1319 -1817 -1314
rect -4299 -1363 -4297 -1358
rect -2113 -1332 -2111 -1327
rect -2103 -1332 -2101 -1327
rect -1775 -1330 -1773 -1320
rect -1767 -1330 -1765 -1320
rect -1733 -1330 -1731 -1320
rect -1725 -1330 -1723 -1320
rect -1688 -1328 -1686 -1323
rect -2731 -1349 -2729 -1344
rect -4255 -1374 -4253 -1364
rect -4247 -1374 -4245 -1364
rect -4213 -1374 -4211 -1364
rect -4205 -1374 -4203 -1364
rect -2781 -1357 -2779 -1352
rect -2771 -1357 -2769 -1352
rect -4168 -1372 -4166 -1367
rect -2615 -1388 -2613 -1383
rect -2665 -1396 -2663 -1391
rect -2655 -1396 -2653 -1391
rect -2424 -1403 -2422 -1393
rect -2414 -1403 -2412 -1393
rect -2375 -1397 -2373 -1392
rect -2914 -1419 -2912 -1409
rect -2904 -1419 -2902 -1409
rect -2865 -1413 -2863 -1408
rect -3485 -1430 -3483 -1420
rect -3475 -1430 -3473 -1420
rect -3436 -1424 -3434 -1419
rect -2727 -1451 -2725 -1446
rect -2240 -1448 -2238 -1443
rect -2777 -1459 -2775 -1454
rect -2767 -1459 -2765 -1454
rect -2290 -1456 -2288 -1451
rect -2280 -1456 -2278 -1451
rect -3194 -1482 -3192 -1477
rect -3309 -1492 -3307 -1487
rect -3244 -1490 -3242 -1485
rect -3234 -1490 -3232 -1485
rect -3359 -1500 -3357 -1495
rect -3349 -1500 -3347 -1495
rect -3819 -1548 -3817 -1538
rect -3809 -1548 -3807 -1538
rect -3770 -1542 -3768 -1537
rect -2910 -1516 -2908 -1506
rect -2900 -1516 -2898 -1506
rect -2861 -1510 -2859 -1505
rect -3665 -1540 -3663 -1535
rect -3480 -1539 -3478 -1529
rect -3470 -1539 -3468 -1529
rect -3431 -1533 -3429 -1528
rect -2425 -1531 -2423 -1521
rect -2415 -1531 -2413 -1521
rect -2376 -1525 -2374 -1520
rect -3715 -1548 -3713 -1543
rect -3705 -1548 -3703 -1543
rect -3815 -1642 -3813 -1637
rect -3770 -1641 -3768 -1631
rect -3760 -1641 -3758 -1631
rect -3721 -1635 -3719 -1630
rect -4265 -1674 -4263 -1669
rect -3463 -1640 -3461 -1635
rect -3418 -1639 -3416 -1629
rect -3408 -1639 -3406 -1629
rect -3369 -1633 -3367 -1628
rect -2227 -1621 -2225 -1616
rect -2182 -1620 -2180 -1610
rect -2172 -1620 -2170 -1610
rect -2133 -1614 -2131 -1609
rect -4221 -1685 -4219 -1675
rect -4213 -1685 -4211 -1675
rect -4179 -1685 -4177 -1675
rect -4171 -1685 -4169 -1675
rect -4134 -1683 -4132 -1678
rect -3815 -1698 -3813 -1693
rect -2902 -1640 -2900 -1635
rect -2857 -1639 -2855 -1629
rect -2847 -1639 -2845 -1629
rect -2808 -1633 -2806 -1628
rect -3612 -1675 -3610 -1670
rect -3662 -1683 -3660 -1678
rect -3652 -1683 -3650 -1678
rect -3463 -1696 -3461 -1691
rect -3260 -1673 -3258 -1668
rect -3310 -1681 -3308 -1676
rect -3300 -1681 -3298 -1676
rect -3768 -1707 -3766 -1697
rect -3758 -1707 -3756 -1697
rect -3719 -1701 -3717 -1696
rect -3416 -1705 -3414 -1695
rect -3406 -1705 -3404 -1695
rect -3367 -1699 -3365 -1694
rect -2902 -1696 -2900 -1691
rect -2699 -1673 -2697 -1668
rect -2749 -1681 -2747 -1676
rect -2739 -1681 -2737 -1676
rect -2227 -1677 -2225 -1672
rect -2024 -1654 -2022 -1649
rect -2074 -1662 -2072 -1657
rect -2064 -1662 -2062 -1657
rect -2180 -1686 -2178 -1676
rect -2170 -1686 -2168 -1676
rect -2131 -1680 -2129 -1675
rect -2855 -1705 -2853 -1695
rect -2845 -1705 -2843 -1695
rect -2806 -1699 -2804 -1694
rect -2193 -1765 -2191 -1755
rect -2183 -1765 -2181 -1755
rect -2144 -1759 -2142 -1754
rect -3413 -1796 -3411 -1786
rect -3403 -1796 -3401 -1786
rect -3364 -1790 -3362 -1785
rect -2863 -1795 -2861 -1785
rect -2853 -1795 -2851 -1785
rect -2814 -1789 -2812 -1784
rect -3800 -1816 -3798 -1806
rect -3790 -1816 -3788 -1806
rect -3751 -1810 -3749 -1805
rect -4246 -1865 -4244 -1860
rect -4202 -1876 -4200 -1866
rect -4194 -1876 -4192 -1866
rect -4160 -1876 -4158 -1866
rect -4152 -1876 -4150 -1866
rect -2947 -1868 -2945 -1863
rect -4115 -1874 -4113 -1869
rect -2903 -1879 -2901 -1869
rect -2895 -1879 -2893 -1869
rect -2861 -1879 -2859 -1869
rect -2853 -1879 -2851 -1869
rect -2709 -1864 -2707 -1859
rect -2260 -1853 -2258 -1848
rect -2816 -1877 -2814 -1872
rect -2665 -1875 -2663 -1865
rect -2657 -1875 -2655 -1865
rect -2623 -1875 -2621 -1865
rect -2615 -1875 -2613 -1865
rect -2216 -1864 -2214 -1854
rect -2208 -1864 -2206 -1854
rect -2174 -1864 -2172 -1854
rect -2166 -1864 -2164 -1854
rect -1943 -1846 -1941 -1841
rect -1899 -1857 -1897 -1847
rect -1891 -1857 -1889 -1847
rect -1857 -1857 -1855 -1847
rect -1849 -1857 -1847 -1847
rect -1812 -1855 -1810 -1850
rect -2129 -1862 -2127 -1857
rect -2578 -1873 -2576 -1868
rect -3622 -2026 -3620 -2021
rect -3578 -2037 -3576 -2027
rect -3570 -2037 -3568 -2027
rect -3536 -2037 -3534 -2027
rect -3528 -2037 -3526 -2027
rect -3323 -2017 -3321 -2012
rect -3279 -2028 -3277 -2018
rect -3271 -2028 -3269 -2018
rect -3237 -2028 -3235 -2018
rect -3229 -2028 -3227 -2018
rect -3192 -2026 -3190 -2021
rect -3491 -2035 -3489 -2030
<< ptransistor >>
rect -3286 -550 -3284 -530
rect -3278 -550 -3276 -530
rect -3234 -550 -3232 -540
rect -3200 -543 -3198 -533
rect -2287 -541 -2285 -521
rect -2279 -541 -2277 -521
rect -1657 -520 -1655 -500
rect -1649 -520 -1647 -500
rect -1605 -520 -1603 -510
rect -1571 -513 -1569 -503
rect -2235 -541 -2233 -531
rect -2201 -534 -2199 -524
rect -3846 -591 -3844 -571
rect -3838 -591 -3836 -571
rect -3794 -591 -3792 -581
rect -3760 -584 -3758 -574
rect -3155 -563 -3153 -553
rect -2156 -554 -2154 -544
rect -1526 -533 -1524 -523
rect -3715 -604 -3713 -594
rect -1880 -732 -1878 -722
rect -1870 -732 -1868 -722
rect -2502 -750 -2500 -740
rect -2492 -750 -2490 -740
rect -1925 -742 -1923 -732
rect -2547 -760 -2545 -750
rect -3223 -776 -3221 -766
rect -3213 -776 -3211 -766
rect -3268 -786 -3266 -776
rect -3174 -779 -3172 -769
rect -2453 -753 -2451 -743
rect -1831 -735 -1829 -725
rect -2394 -796 -2392 -776
rect -2384 -796 -2382 -776
rect -1772 -778 -1770 -758
rect -1762 -778 -1760 -758
rect -1722 -775 -1720 -765
rect -2344 -793 -2342 -783
rect -3115 -822 -3113 -802
rect -3105 -822 -3103 -802
rect -3065 -819 -3063 -809
rect -2547 -816 -2545 -806
rect -2500 -816 -2498 -806
rect -2490 -816 -2488 -806
rect -3268 -842 -3266 -832
rect -3221 -842 -3219 -832
rect -3211 -842 -3209 -832
rect -3172 -845 -3170 -835
rect -2451 -819 -2449 -809
rect -1925 -798 -1923 -788
rect -1878 -798 -1876 -788
rect -1868 -798 -1866 -788
rect -1829 -801 -1827 -791
rect -3768 -1022 -3766 -1012
rect -3758 -1022 -3756 -1012
rect -3813 -1032 -3811 -1022
rect -3719 -1025 -3717 -1015
rect -3660 -1068 -3658 -1048
rect -3650 -1068 -3648 -1048
rect -3610 -1065 -3608 -1055
rect -3813 -1088 -3811 -1078
rect -3766 -1088 -3764 -1078
rect -3756 -1088 -3754 -1078
rect -3717 -1091 -3715 -1081
rect -2428 -1128 -2426 -1118
rect -2418 -1128 -2416 -1118
rect -2379 -1131 -2377 -1121
rect -2289 -1187 -2287 -1167
rect -2279 -1187 -2277 -1167
rect -2239 -1184 -2237 -1174
rect -2429 -1251 -2427 -1241
rect -2419 -1251 -2417 -1241
rect -2380 -1254 -2378 -1244
rect -2913 -1284 -2911 -1274
rect -2903 -1284 -2901 -1274
rect -2864 -1287 -2862 -1277
rect -2113 -1307 -2111 -1287
rect -2103 -1307 -2101 -1287
rect -2063 -1304 -2061 -1294
rect -1928 -1298 -1926 -1278
rect -1918 -1298 -1916 -1278
rect -1878 -1295 -1876 -1285
rect -1819 -1295 -1817 -1275
rect -1811 -1295 -1809 -1275
rect -1767 -1295 -1765 -1285
rect -1733 -1288 -1731 -1278
rect -4299 -1339 -4297 -1319
rect -4291 -1339 -4289 -1319
rect -4247 -1339 -4245 -1329
rect -4213 -1332 -4211 -1322
rect -2781 -1332 -2779 -1312
rect -2771 -1332 -2769 -1312
rect -2731 -1329 -2729 -1319
rect -1688 -1308 -1686 -1298
rect -4168 -1352 -4166 -1342
rect -2665 -1371 -2663 -1351
rect -2655 -1371 -2653 -1351
rect -2615 -1368 -2613 -1358
rect -2914 -1390 -2912 -1380
rect -2904 -1390 -2902 -1380
rect -3485 -1401 -3483 -1391
rect -3475 -1401 -3473 -1391
rect -3436 -1404 -3434 -1394
rect -2865 -1393 -2863 -1383
rect -2424 -1374 -2422 -1364
rect -2414 -1374 -2412 -1364
rect -2375 -1377 -2373 -1367
rect -2777 -1434 -2775 -1414
rect -2767 -1434 -2765 -1414
rect -2727 -1431 -2725 -1421
rect -2290 -1431 -2288 -1411
rect -2280 -1431 -2278 -1411
rect -2240 -1428 -2238 -1418
rect -3359 -1475 -3357 -1455
rect -3349 -1475 -3347 -1455
rect -3309 -1472 -3307 -1462
rect -3244 -1465 -3242 -1445
rect -3234 -1465 -3232 -1445
rect -3194 -1462 -3192 -1452
rect -2910 -1487 -2908 -1477
rect -2900 -1487 -2898 -1477
rect -3819 -1519 -3817 -1509
rect -3809 -1519 -3807 -1509
rect -3770 -1522 -3768 -1512
rect -3715 -1523 -3713 -1503
rect -3705 -1523 -3703 -1503
rect -3480 -1510 -3478 -1500
rect -3470 -1510 -3468 -1500
rect -3665 -1520 -3663 -1510
rect -3431 -1513 -3429 -1503
rect -2861 -1490 -2859 -1480
rect -2425 -1502 -2423 -1492
rect -2415 -1502 -2413 -1492
rect -2376 -1505 -2374 -1495
rect -2182 -1591 -2180 -1581
rect -2172 -1591 -2170 -1581
rect -3770 -1612 -3768 -1602
rect -3760 -1612 -3758 -1602
rect -3815 -1622 -3813 -1612
rect -4265 -1650 -4263 -1630
rect -4257 -1650 -4255 -1630
rect -4213 -1650 -4211 -1640
rect -4179 -1643 -4177 -1633
rect -3721 -1615 -3719 -1605
rect -3418 -1610 -3416 -1600
rect -3408 -1610 -3406 -1600
rect -3463 -1620 -3461 -1610
rect -3369 -1613 -3367 -1603
rect -2857 -1610 -2855 -1600
rect -2847 -1610 -2845 -1600
rect -2227 -1601 -2225 -1591
rect -2902 -1620 -2900 -1610
rect -4134 -1663 -4132 -1653
rect -3662 -1658 -3660 -1638
rect -3652 -1658 -3650 -1638
rect -2808 -1613 -2806 -1603
rect -2133 -1594 -2131 -1584
rect -3612 -1655 -3610 -1645
rect -3815 -1678 -3813 -1668
rect -3768 -1678 -3766 -1668
rect -3758 -1678 -3756 -1668
rect -3719 -1681 -3717 -1671
rect -3310 -1656 -3308 -1636
rect -3300 -1656 -3298 -1636
rect -3260 -1653 -3258 -1643
rect -3463 -1676 -3461 -1666
rect -3416 -1676 -3414 -1666
rect -3406 -1676 -3404 -1666
rect -3367 -1679 -3365 -1669
rect -2749 -1656 -2747 -1636
rect -2739 -1656 -2737 -1636
rect -2074 -1637 -2072 -1617
rect -2064 -1637 -2062 -1617
rect -2024 -1634 -2022 -1624
rect -2699 -1653 -2697 -1643
rect -2902 -1676 -2900 -1666
rect -2855 -1676 -2853 -1666
rect -2845 -1676 -2843 -1666
rect -2806 -1679 -2804 -1669
rect -2227 -1657 -2225 -1647
rect -2180 -1657 -2178 -1647
rect -2170 -1657 -2168 -1647
rect -2131 -1660 -2129 -1650
rect -2193 -1736 -2191 -1726
rect -2183 -1736 -2181 -1726
rect -2144 -1739 -2142 -1729
rect -3413 -1767 -3411 -1757
rect -3403 -1767 -3401 -1757
rect -3800 -1787 -3798 -1777
rect -3790 -1787 -3788 -1777
rect -3751 -1790 -3749 -1780
rect -3364 -1770 -3362 -1760
rect -2863 -1766 -2861 -1756
rect -2853 -1766 -2851 -1756
rect -2814 -1769 -2812 -1759
rect -4246 -1841 -4244 -1821
rect -4238 -1841 -4236 -1821
rect -4194 -1841 -4192 -1831
rect -4160 -1834 -4158 -1824
rect -2947 -1844 -2945 -1824
rect -2939 -1844 -2937 -1824
rect -2895 -1844 -2893 -1834
rect -2861 -1837 -2859 -1827
rect -4115 -1854 -4113 -1844
rect -2709 -1840 -2707 -1820
rect -2701 -1840 -2699 -1820
rect -2657 -1840 -2655 -1830
rect -2623 -1833 -2621 -1823
rect -2260 -1829 -2258 -1809
rect -2252 -1829 -2250 -1809
rect -2208 -1829 -2206 -1819
rect -2174 -1822 -2172 -1812
rect -1943 -1822 -1941 -1802
rect -1935 -1822 -1933 -1802
rect -1891 -1822 -1889 -1812
rect -1857 -1815 -1855 -1805
rect -2816 -1857 -2814 -1847
rect -2578 -1853 -2576 -1843
rect -2129 -1842 -2127 -1832
rect -1812 -1835 -1810 -1825
rect -3622 -2002 -3620 -1982
rect -3614 -2002 -3612 -1982
rect -3570 -2002 -3568 -1992
rect -3536 -1995 -3534 -1985
rect -3323 -1993 -3321 -1973
rect -3315 -1993 -3313 -1973
rect -3271 -1993 -3269 -1983
rect -3237 -1986 -3235 -1976
rect -3491 -2015 -3489 -2005
rect -3192 -2006 -3190 -1996
<< ndiffusion >>
rect -3287 -574 -3286 -569
rect -3284 -574 -3275 -569
rect -3847 -615 -3846 -610
rect -3844 -615 -3835 -610
rect -3243 -585 -3242 -575
rect -3240 -585 -3234 -575
rect -3232 -585 -3224 -575
rect -3201 -585 -3200 -575
rect -3198 -585 -3192 -575
rect -3190 -585 -3189 -575
rect -2288 -565 -2287 -560
rect -2285 -565 -2276 -560
rect -1658 -544 -1657 -539
rect -1655 -544 -1646 -539
rect -2244 -576 -2243 -566
rect -2241 -576 -2235 -566
rect -2233 -576 -2225 -566
rect -2202 -576 -2201 -566
rect -2199 -576 -2193 -566
rect -2191 -576 -2190 -566
rect -1614 -555 -1613 -545
rect -1611 -555 -1605 -545
rect -1603 -555 -1595 -545
rect -1572 -555 -1571 -545
rect -1569 -555 -1563 -545
rect -1561 -555 -1560 -545
rect -1528 -553 -1526 -548
rect -1524 -553 -1514 -548
rect -2158 -574 -2156 -569
rect -2154 -574 -2144 -569
rect -3157 -583 -3155 -578
rect -3153 -583 -3143 -578
rect -3803 -626 -3802 -616
rect -3800 -626 -3794 -616
rect -3792 -626 -3784 -616
rect -3761 -626 -3760 -616
rect -3758 -626 -3752 -616
rect -3750 -626 -3749 -616
rect -3717 -624 -3715 -619
rect -3713 -624 -3703 -619
rect -1927 -762 -1925 -757
rect -1923 -762 -1913 -757
rect -1881 -761 -1880 -751
rect -1878 -761 -1870 -751
rect -1868 -761 -1867 -751
rect -1833 -755 -1831 -750
rect -1829 -755 -1819 -750
rect -2549 -780 -2547 -775
rect -2545 -780 -2535 -775
rect -2503 -779 -2502 -769
rect -2500 -779 -2492 -769
rect -2490 -779 -2489 -769
rect -2455 -773 -2453 -768
rect -2451 -773 -2441 -768
rect -3270 -806 -3268 -801
rect -3266 -806 -3256 -801
rect -3224 -805 -3223 -795
rect -3221 -805 -3213 -795
rect -3211 -805 -3210 -795
rect -3176 -799 -3174 -794
rect -3172 -799 -3162 -794
rect -3270 -862 -3268 -857
rect -3266 -862 -3256 -857
rect -3067 -839 -3065 -834
rect -3063 -839 -3053 -834
rect -2549 -836 -2547 -831
rect -2545 -836 -2535 -831
rect -2346 -813 -2344 -808
rect -2342 -813 -2332 -808
rect -2395 -821 -2394 -816
rect -2392 -821 -2391 -816
rect -2385 -821 -2384 -816
rect -2382 -821 -2381 -816
rect -1927 -818 -1925 -813
rect -1923 -818 -1913 -813
rect -1724 -795 -1722 -790
rect -1720 -795 -1710 -790
rect -1773 -803 -1772 -798
rect -1770 -803 -1769 -798
rect -1763 -803 -1762 -798
rect -1760 -803 -1759 -798
rect -1879 -827 -1878 -817
rect -1876 -827 -1868 -817
rect -1866 -827 -1865 -817
rect -1831 -821 -1829 -816
rect -1827 -821 -1817 -816
rect -3116 -847 -3115 -842
rect -3113 -847 -3112 -842
rect -3106 -847 -3105 -842
rect -3103 -847 -3102 -842
rect -2501 -845 -2500 -835
rect -2498 -845 -2490 -835
rect -2488 -845 -2487 -835
rect -2453 -839 -2451 -834
rect -2449 -839 -2439 -834
rect -3222 -871 -3221 -861
rect -3219 -871 -3211 -861
rect -3209 -871 -3208 -861
rect -3174 -865 -3172 -860
rect -3170 -865 -3160 -860
rect -3815 -1052 -3813 -1047
rect -3811 -1052 -3801 -1047
rect -3769 -1051 -3768 -1041
rect -3766 -1051 -3758 -1041
rect -3756 -1051 -3755 -1041
rect -3721 -1045 -3719 -1040
rect -3717 -1045 -3707 -1040
rect -3815 -1108 -3813 -1103
rect -3811 -1108 -3801 -1103
rect -3612 -1085 -3610 -1080
rect -3608 -1085 -3598 -1080
rect -3661 -1093 -3660 -1088
rect -3658 -1093 -3657 -1088
rect -3651 -1093 -3650 -1088
rect -3648 -1093 -3647 -1088
rect -3767 -1117 -3766 -1107
rect -3764 -1117 -3756 -1107
rect -3754 -1117 -3753 -1107
rect -3719 -1111 -3717 -1106
rect -3715 -1111 -3705 -1106
rect -2429 -1157 -2428 -1147
rect -2426 -1157 -2418 -1147
rect -2416 -1157 -2415 -1147
rect -2381 -1151 -2379 -1146
rect -2377 -1151 -2367 -1146
rect -2241 -1204 -2239 -1199
rect -2237 -1204 -2227 -1199
rect -2290 -1212 -2289 -1207
rect -2287 -1212 -2286 -1207
rect -2280 -1212 -2279 -1207
rect -2277 -1212 -2276 -1207
rect -2430 -1280 -2429 -1270
rect -2427 -1280 -2419 -1270
rect -2417 -1280 -2416 -1270
rect -2382 -1274 -2380 -1269
rect -2378 -1274 -2368 -1269
rect -2914 -1313 -2913 -1303
rect -2911 -1313 -2903 -1303
rect -2901 -1313 -2900 -1303
rect -2866 -1307 -2864 -1302
rect -2862 -1307 -2852 -1302
rect -1880 -1315 -1878 -1310
rect -1876 -1315 -1866 -1310
rect -2065 -1324 -2063 -1319
rect -2061 -1324 -2051 -1319
rect -1929 -1323 -1928 -1318
rect -1926 -1323 -1925 -1318
rect -1919 -1323 -1918 -1318
rect -1916 -1323 -1915 -1318
rect -1820 -1319 -1819 -1314
rect -1817 -1319 -1808 -1314
rect -4300 -1363 -4299 -1358
rect -4297 -1363 -4288 -1358
rect -2114 -1332 -2113 -1327
rect -2111 -1332 -2110 -1327
rect -2104 -1332 -2103 -1327
rect -2101 -1332 -2100 -1327
rect -1776 -1330 -1775 -1320
rect -1773 -1330 -1767 -1320
rect -1765 -1330 -1757 -1320
rect -1734 -1330 -1733 -1320
rect -1731 -1330 -1725 -1320
rect -1723 -1330 -1722 -1320
rect -1690 -1328 -1688 -1323
rect -1686 -1328 -1676 -1323
rect -2733 -1349 -2731 -1344
rect -2729 -1349 -2719 -1344
rect -4256 -1374 -4255 -1364
rect -4253 -1374 -4247 -1364
rect -4245 -1374 -4237 -1364
rect -4214 -1374 -4213 -1364
rect -4211 -1374 -4205 -1364
rect -4203 -1374 -4202 -1364
rect -2782 -1357 -2781 -1352
rect -2779 -1357 -2778 -1352
rect -2772 -1357 -2771 -1352
rect -2769 -1357 -2768 -1352
rect -4170 -1372 -4168 -1367
rect -4166 -1372 -4156 -1367
rect -2617 -1388 -2615 -1383
rect -2613 -1388 -2603 -1383
rect -2666 -1396 -2665 -1391
rect -2663 -1396 -2662 -1391
rect -2656 -1396 -2655 -1391
rect -2653 -1396 -2652 -1391
rect -2425 -1403 -2424 -1393
rect -2422 -1403 -2414 -1393
rect -2412 -1403 -2411 -1393
rect -2377 -1397 -2375 -1392
rect -2373 -1397 -2363 -1392
rect -2915 -1419 -2914 -1409
rect -2912 -1419 -2904 -1409
rect -2902 -1419 -2901 -1409
rect -2867 -1413 -2865 -1408
rect -2863 -1413 -2853 -1408
rect -3486 -1430 -3485 -1420
rect -3483 -1430 -3475 -1420
rect -3473 -1430 -3472 -1420
rect -3438 -1424 -3436 -1419
rect -3434 -1424 -3424 -1419
rect -2729 -1451 -2727 -1446
rect -2725 -1451 -2715 -1446
rect -2242 -1448 -2240 -1443
rect -2238 -1448 -2228 -1443
rect -2778 -1459 -2777 -1454
rect -2775 -1459 -2774 -1454
rect -2768 -1459 -2767 -1454
rect -2765 -1459 -2764 -1454
rect -2291 -1456 -2290 -1451
rect -2288 -1456 -2287 -1451
rect -2281 -1456 -2280 -1451
rect -2278 -1456 -2277 -1451
rect -3196 -1482 -3194 -1477
rect -3192 -1482 -3182 -1477
rect -3311 -1492 -3309 -1487
rect -3307 -1492 -3297 -1487
rect -3245 -1490 -3244 -1485
rect -3242 -1490 -3241 -1485
rect -3235 -1490 -3234 -1485
rect -3232 -1490 -3231 -1485
rect -3360 -1500 -3359 -1495
rect -3357 -1500 -3356 -1495
rect -3350 -1500 -3349 -1495
rect -3347 -1500 -3346 -1495
rect -3820 -1548 -3819 -1538
rect -3817 -1548 -3809 -1538
rect -3807 -1548 -3806 -1538
rect -3772 -1542 -3770 -1537
rect -3768 -1542 -3758 -1537
rect -2911 -1516 -2910 -1506
rect -2908 -1516 -2900 -1506
rect -2898 -1516 -2897 -1506
rect -2863 -1510 -2861 -1505
rect -2859 -1510 -2849 -1505
rect -3667 -1540 -3665 -1535
rect -3663 -1540 -3653 -1535
rect -3481 -1539 -3480 -1529
rect -3478 -1539 -3470 -1529
rect -3468 -1539 -3467 -1529
rect -3433 -1533 -3431 -1528
rect -3429 -1533 -3419 -1528
rect -2426 -1531 -2425 -1521
rect -2423 -1531 -2415 -1521
rect -2413 -1531 -2412 -1521
rect -2378 -1525 -2376 -1520
rect -2374 -1525 -2364 -1520
rect -3716 -1548 -3715 -1543
rect -3713 -1548 -3712 -1543
rect -3706 -1548 -3705 -1543
rect -3703 -1548 -3702 -1543
rect -3817 -1642 -3815 -1637
rect -3813 -1642 -3803 -1637
rect -3771 -1641 -3770 -1631
rect -3768 -1641 -3760 -1631
rect -3758 -1641 -3757 -1631
rect -3723 -1635 -3721 -1630
rect -3719 -1635 -3709 -1630
rect -4266 -1674 -4265 -1669
rect -4263 -1674 -4254 -1669
rect -3465 -1640 -3463 -1635
rect -3461 -1640 -3451 -1635
rect -3419 -1639 -3418 -1629
rect -3416 -1639 -3408 -1629
rect -3406 -1639 -3405 -1629
rect -3371 -1633 -3369 -1628
rect -3367 -1633 -3357 -1628
rect -2229 -1621 -2227 -1616
rect -2225 -1621 -2215 -1616
rect -2183 -1620 -2182 -1610
rect -2180 -1620 -2172 -1610
rect -2170 -1620 -2169 -1610
rect -2135 -1614 -2133 -1609
rect -2131 -1614 -2121 -1609
rect -4222 -1685 -4221 -1675
rect -4219 -1685 -4213 -1675
rect -4211 -1685 -4203 -1675
rect -4180 -1685 -4179 -1675
rect -4177 -1685 -4171 -1675
rect -4169 -1685 -4168 -1675
rect -4136 -1683 -4134 -1678
rect -4132 -1683 -4122 -1678
rect -3817 -1698 -3815 -1693
rect -3813 -1698 -3803 -1693
rect -2904 -1640 -2902 -1635
rect -2900 -1640 -2890 -1635
rect -2858 -1639 -2857 -1629
rect -2855 -1639 -2847 -1629
rect -2845 -1639 -2844 -1629
rect -2810 -1633 -2808 -1628
rect -2806 -1633 -2796 -1628
rect -3614 -1675 -3612 -1670
rect -3610 -1675 -3600 -1670
rect -3663 -1683 -3662 -1678
rect -3660 -1683 -3659 -1678
rect -3653 -1683 -3652 -1678
rect -3650 -1683 -3649 -1678
rect -3465 -1696 -3463 -1691
rect -3461 -1696 -3451 -1691
rect -3262 -1673 -3260 -1668
rect -3258 -1673 -3248 -1668
rect -3311 -1681 -3310 -1676
rect -3308 -1681 -3307 -1676
rect -3301 -1681 -3300 -1676
rect -3298 -1681 -3297 -1676
rect -3769 -1707 -3768 -1697
rect -3766 -1707 -3758 -1697
rect -3756 -1707 -3755 -1697
rect -3721 -1701 -3719 -1696
rect -3717 -1701 -3707 -1696
rect -3417 -1705 -3416 -1695
rect -3414 -1705 -3406 -1695
rect -3404 -1705 -3403 -1695
rect -3369 -1699 -3367 -1694
rect -3365 -1699 -3355 -1694
rect -2904 -1696 -2902 -1691
rect -2900 -1696 -2890 -1691
rect -2701 -1673 -2699 -1668
rect -2697 -1673 -2687 -1668
rect -2750 -1681 -2749 -1676
rect -2747 -1681 -2746 -1676
rect -2740 -1681 -2739 -1676
rect -2737 -1681 -2736 -1676
rect -2229 -1677 -2227 -1672
rect -2225 -1677 -2215 -1672
rect -2026 -1654 -2024 -1649
rect -2022 -1654 -2012 -1649
rect -2075 -1662 -2074 -1657
rect -2072 -1662 -2071 -1657
rect -2065 -1662 -2064 -1657
rect -2062 -1662 -2061 -1657
rect -2181 -1686 -2180 -1676
rect -2178 -1686 -2170 -1676
rect -2168 -1686 -2167 -1676
rect -2133 -1680 -2131 -1675
rect -2129 -1680 -2119 -1675
rect -2856 -1705 -2855 -1695
rect -2853 -1705 -2845 -1695
rect -2843 -1705 -2842 -1695
rect -2808 -1699 -2806 -1694
rect -2804 -1699 -2794 -1694
rect -2194 -1765 -2193 -1755
rect -2191 -1765 -2183 -1755
rect -2181 -1765 -2180 -1755
rect -2146 -1759 -2144 -1754
rect -2142 -1759 -2132 -1754
rect -3414 -1796 -3413 -1786
rect -3411 -1796 -3403 -1786
rect -3401 -1796 -3400 -1786
rect -3366 -1790 -3364 -1785
rect -3362 -1790 -3352 -1785
rect -2864 -1795 -2863 -1785
rect -2861 -1795 -2853 -1785
rect -2851 -1795 -2850 -1785
rect -2816 -1789 -2814 -1784
rect -2812 -1789 -2802 -1784
rect -3801 -1816 -3800 -1806
rect -3798 -1816 -3790 -1806
rect -3788 -1816 -3787 -1806
rect -3753 -1810 -3751 -1805
rect -3749 -1810 -3739 -1805
rect -4247 -1865 -4246 -1860
rect -4244 -1865 -4235 -1860
rect -4203 -1876 -4202 -1866
rect -4200 -1876 -4194 -1866
rect -4192 -1876 -4184 -1866
rect -4161 -1876 -4160 -1866
rect -4158 -1876 -4152 -1866
rect -4150 -1876 -4149 -1866
rect -2948 -1868 -2947 -1863
rect -2945 -1868 -2936 -1863
rect -4117 -1874 -4115 -1869
rect -4113 -1874 -4103 -1869
rect -2904 -1879 -2903 -1869
rect -2901 -1879 -2895 -1869
rect -2893 -1879 -2885 -1869
rect -2862 -1879 -2861 -1869
rect -2859 -1879 -2853 -1869
rect -2851 -1879 -2850 -1869
rect -2710 -1864 -2709 -1859
rect -2707 -1864 -2698 -1859
rect -2261 -1853 -2260 -1848
rect -2258 -1853 -2249 -1848
rect -2818 -1877 -2816 -1872
rect -2814 -1877 -2804 -1872
rect -2666 -1875 -2665 -1865
rect -2663 -1875 -2657 -1865
rect -2655 -1875 -2647 -1865
rect -2624 -1875 -2623 -1865
rect -2621 -1875 -2615 -1865
rect -2613 -1875 -2612 -1865
rect -2217 -1864 -2216 -1854
rect -2214 -1864 -2208 -1854
rect -2206 -1864 -2198 -1854
rect -2175 -1864 -2174 -1854
rect -2172 -1864 -2166 -1854
rect -2164 -1864 -2163 -1854
rect -1944 -1846 -1943 -1841
rect -1941 -1846 -1932 -1841
rect -1900 -1857 -1899 -1847
rect -1897 -1857 -1891 -1847
rect -1889 -1857 -1881 -1847
rect -1858 -1857 -1857 -1847
rect -1855 -1857 -1849 -1847
rect -1847 -1857 -1846 -1847
rect -1814 -1855 -1812 -1850
rect -1810 -1855 -1800 -1850
rect -2131 -1862 -2129 -1857
rect -2127 -1862 -2117 -1857
rect -2580 -1873 -2578 -1868
rect -2576 -1873 -2566 -1868
rect -3623 -2026 -3622 -2021
rect -3620 -2026 -3611 -2021
rect -3579 -2037 -3578 -2027
rect -3576 -2037 -3570 -2027
rect -3568 -2037 -3560 -2027
rect -3537 -2037 -3536 -2027
rect -3534 -2037 -3528 -2027
rect -3526 -2037 -3525 -2027
rect -3324 -2017 -3323 -2012
rect -3321 -2017 -3312 -2012
rect -3280 -2028 -3279 -2018
rect -3277 -2028 -3271 -2018
rect -3269 -2028 -3261 -2018
rect -3238 -2028 -3237 -2018
rect -3235 -2028 -3229 -2018
rect -3227 -2028 -3226 -2018
rect -3194 -2026 -3192 -2021
rect -3190 -2026 -3180 -2021
rect -3493 -2035 -3491 -2030
rect -3489 -2035 -3479 -2030
<< pdiffusion >>
rect -3287 -550 -3286 -530
rect -3284 -550 -3278 -530
rect -3276 -550 -3275 -530
rect -3235 -550 -3234 -540
rect -3232 -550 -3231 -540
rect -3201 -543 -3200 -533
rect -3198 -543 -3197 -533
rect -2288 -541 -2287 -521
rect -2285 -541 -2279 -521
rect -2277 -541 -2276 -521
rect -1658 -520 -1657 -500
rect -1655 -520 -1649 -500
rect -1647 -520 -1646 -500
rect -1606 -520 -1605 -510
rect -1603 -520 -1602 -510
rect -1572 -513 -1571 -503
rect -1569 -513 -1568 -503
rect -2236 -541 -2235 -531
rect -2233 -541 -2232 -531
rect -2202 -534 -2201 -524
rect -2199 -534 -2198 -524
rect -3847 -591 -3846 -571
rect -3844 -591 -3838 -571
rect -3836 -591 -3835 -571
rect -3795 -591 -3794 -581
rect -3792 -591 -3791 -581
rect -3761 -584 -3760 -574
rect -3758 -584 -3757 -574
rect -3157 -563 -3155 -553
rect -3153 -563 -3143 -553
rect -2158 -554 -2156 -544
rect -2154 -554 -2144 -544
rect -1528 -533 -1526 -523
rect -1524 -533 -1514 -523
rect -3717 -604 -3715 -594
rect -3713 -604 -3703 -594
rect -1881 -732 -1880 -722
rect -1878 -732 -1876 -722
rect -1872 -732 -1870 -722
rect -1868 -732 -1867 -722
rect -2503 -750 -2502 -740
rect -2500 -750 -2498 -740
rect -2494 -750 -2492 -740
rect -2490 -750 -2489 -740
rect -1927 -742 -1925 -732
rect -1923 -742 -1913 -732
rect -2549 -760 -2547 -750
rect -2545 -760 -2535 -750
rect -3224 -776 -3223 -766
rect -3221 -776 -3219 -766
rect -3215 -776 -3213 -766
rect -3211 -776 -3210 -766
rect -3270 -786 -3268 -776
rect -3266 -786 -3256 -776
rect -3176 -779 -3174 -769
rect -3172 -779 -3162 -769
rect -2455 -753 -2453 -743
rect -2451 -753 -2441 -743
rect -1833 -735 -1831 -725
rect -1829 -735 -1819 -725
rect -2395 -796 -2394 -776
rect -2392 -796 -2384 -776
rect -2382 -796 -2381 -776
rect -1773 -778 -1772 -758
rect -1770 -778 -1762 -758
rect -1760 -778 -1759 -758
rect -1724 -775 -1722 -765
rect -1720 -775 -1710 -765
rect -2346 -793 -2344 -783
rect -2342 -793 -2332 -783
rect -3116 -822 -3115 -802
rect -3113 -822 -3105 -802
rect -3103 -822 -3102 -802
rect -3067 -819 -3065 -809
rect -3063 -819 -3053 -809
rect -2549 -816 -2547 -806
rect -2545 -816 -2535 -806
rect -2501 -816 -2500 -806
rect -2498 -816 -2496 -806
rect -2492 -816 -2490 -806
rect -2488 -816 -2487 -806
rect -3270 -842 -3268 -832
rect -3266 -842 -3256 -832
rect -3222 -842 -3221 -832
rect -3219 -842 -3217 -832
rect -3213 -842 -3211 -832
rect -3209 -842 -3208 -832
rect -3174 -845 -3172 -835
rect -3170 -845 -3160 -835
rect -2453 -819 -2451 -809
rect -2449 -819 -2439 -809
rect -1927 -798 -1925 -788
rect -1923 -798 -1913 -788
rect -1879 -798 -1878 -788
rect -1876 -798 -1874 -788
rect -1870 -798 -1868 -788
rect -1866 -798 -1865 -788
rect -1831 -801 -1829 -791
rect -1827 -801 -1817 -791
rect -3769 -1022 -3768 -1012
rect -3766 -1022 -3764 -1012
rect -3760 -1022 -3758 -1012
rect -3756 -1022 -3755 -1012
rect -3815 -1032 -3813 -1022
rect -3811 -1032 -3801 -1022
rect -3721 -1025 -3719 -1015
rect -3717 -1025 -3707 -1015
rect -3661 -1068 -3660 -1048
rect -3658 -1068 -3650 -1048
rect -3648 -1068 -3647 -1048
rect -3612 -1065 -3610 -1055
rect -3608 -1065 -3598 -1055
rect -3815 -1088 -3813 -1078
rect -3811 -1088 -3801 -1078
rect -3767 -1088 -3766 -1078
rect -3764 -1088 -3762 -1078
rect -3758 -1088 -3756 -1078
rect -3754 -1088 -3753 -1078
rect -3719 -1091 -3717 -1081
rect -3715 -1091 -3705 -1081
rect -2429 -1128 -2428 -1118
rect -2426 -1128 -2424 -1118
rect -2420 -1128 -2418 -1118
rect -2416 -1128 -2415 -1118
rect -2381 -1131 -2379 -1121
rect -2377 -1131 -2367 -1121
rect -2290 -1187 -2289 -1167
rect -2287 -1187 -2279 -1167
rect -2277 -1187 -2276 -1167
rect -2241 -1184 -2239 -1174
rect -2237 -1184 -2227 -1174
rect -2430 -1251 -2429 -1241
rect -2427 -1251 -2425 -1241
rect -2421 -1251 -2419 -1241
rect -2417 -1251 -2416 -1241
rect -2382 -1254 -2380 -1244
rect -2378 -1254 -2368 -1244
rect -2914 -1284 -2913 -1274
rect -2911 -1284 -2909 -1274
rect -2905 -1284 -2903 -1274
rect -2901 -1284 -2900 -1274
rect -2866 -1287 -2864 -1277
rect -2862 -1287 -2852 -1277
rect -2114 -1307 -2113 -1287
rect -2111 -1307 -2103 -1287
rect -2101 -1307 -2100 -1287
rect -2065 -1304 -2063 -1294
rect -2061 -1304 -2051 -1294
rect -1929 -1298 -1928 -1278
rect -1926 -1298 -1918 -1278
rect -1916 -1298 -1915 -1278
rect -1880 -1295 -1878 -1285
rect -1876 -1295 -1866 -1285
rect -1820 -1295 -1819 -1275
rect -1817 -1295 -1811 -1275
rect -1809 -1295 -1808 -1275
rect -1768 -1295 -1767 -1285
rect -1765 -1295 -1764 -1285
rect -1734 -1288 -1733 -1278
rect -1731 -1288 -1730 -1278
rect -4300 -1339 -4299 -1319
rect -4297 -1339 -4291 -1319
rect -4289 -1339 -4288 -1319
rect -4248 -1339 -4247 -1329
rect -4245 -1339 -4244 -1329
rect -4214 -1332 -4213 -1322
rect -4211 -1332 -4210 -1322
rect -2782 -1332 -2781 -1312
rect -2779 -1332 -2771 -1312
rect -2769 -1332 -2768 -1312
rect -2733 -1329 -2731 -1319
rect -2729 -1329 -2719 -1319
rect -1690 -1308 -1688 -1298
rect -1686 -1308 -1676 -1298
rect -4170 -1352 -4168 -1342
rect -4166 -1352 -4156 -1342
rect -2666 -1371 -2665 -1351
rect -2663 -1371 -2655 -1351
rect -2653 -1371 -2652 -1351
rect -2617 -1368 -2615 -1358
rect -2613 -1368 -2603 -1358
rect -2915 -1390 -2914 -1380
rect -2912 -1390 -2910 -1380
rect -2906 -1390 -2904 -1380
rect -2902 -1390 -2901 -1380
rect -3486 -1401 -3485 -1391
rect -3483 -1401 -3481 -1391
rect -3477 -1401 -3475 -1391
rect -3473 -1401 -3472 -1391
rect -3438 -1404 -3436 -1394
rect -3434 -1404 -3424 -1394
rect -2867 -1393 -2865 -1383
rect -2863 -1393 -2853 -1383
rect -2425 -1374 -2424 -1364
rect -2422 -1374 -2420 -1364
rect -2416 -1374 -2414 -1364
rect -2412 -1374 -2411 -1364
rect -2377 -1377 -2375 -1367
rect -2373 -1377 -2363 -1367
rect -2778 -1434 -2777 -1414
rect -2775 -1434 -2767 -1414
rect -2765 -1434 -2764 -1414
rect -2729 -1431 -2727 -1421
rect -2725 -1431 -2715 -1421
rect -2291 -1431 -2290 -1411
rect -2288 -1431 -2280 -1411
rect -2278 -1431 -2277 -1411
rect -2242 -1428 -2240 -1418
rect -2238 -1428 -2228 -1418
rect -3360 -1475 -3359 -1455
rect -3357 -1475 -3349 -1455
rect -3347 -1475 -3346 -1455
rect -3311 -1472 -3309 -1462
rect -3307 -1472 -3297 -1462
rect -3245 -1465 -3244 -1445
rect -3242 -1465 -3234 -1445
rect -3232 -1465 -3231 -1445
rect -3196 -1462 -3194 -1452
rect -3192 -1462 -3182 -1452
rect -2911 -1487 -2910 -1477
rect -2908 -1487 -2906 -1477
rect -2902 -1487 -2900 -1477
rect -2898 -1487 -2897 -1477
rect -3820 -1519 -3819 -1509
rect -3817 -1519 -3815 -1509
rect -3811 -1519 -3809 -1509
rect -3807 -1519 -3806 -1509
rect -3772 -1522 -3770 -1512
rect -3768 -1522 -3758 -1512
rect -3716 -1523 -3715 -1503
rect -3713 -1523 -3705 -1503
rect -3703 -1523 -3702 -1503
rect -3481 -1510 -3480 -1500
rect -3478 -1510 -3476 -1500
rect -3472 -1510 -3470 -1500
rect -3468 -1510 -3467 -1500
rect -3667 -1520 -3665 -1510
rect -3663 -1520 -3653 -1510
rect -3433 -1513 -3431 -1503
rect -3429 -1513 -3419 -1503
rect -2863 -1490 -2861 -1480
rect -2859 -1490 -2849 -1480
rect -2426 -1502 -2425 -1492
rect -2423 -1502 -2421 -1492
rect -2417 -1502 -2415 -1492
rect -2413 -1502 -2412 -1492
rect -2378 -1505 -2376 -1495
rect -2374 -1505 -2364 -1495
rect -2183 -1591 -2182 -1581
rect -2180 -1591 -2178 -1581
rect -2174 -1591 -2172 -1581
rect -2170 -1591 -2169 -1581
rect -3771 -1612 -3770 -1602
rect -3768 -1612 -3766 -1602
rect -3762 -1612 -3760 -1602
rect -3758 -1612 -3757 -1602
rect -3817 -1622 -3815 -1612
rect -3813 -1622 -3803 -1612
rect -4266 -1650 -4265 -1630
rect -4263 -1650 -4257 -1630
rect -4255 -1650 -4254 -1630
rect -4214 -1650 -4213 -1640
rect -4211 -1650 -4210 -1640
rect -4180 -1643 -4179 -1633
rect -4177 -1643 -4176 -1633
rect -3723 -1615 -3721 -1605
rect -3719 -1615 -3709 -1605
rect -3419 -1610 -3418 -1600
rect -3416 -1610 -3414 -1600
rect -3410 -1610 -3408 -1600
rect -3406 -1610 -3405 -1600
rect -3465 -1620 -3463 -1610
rect -3461 -1620 -3451 -1610
rect -3371 -1613 -3369 -1603
rect -3367 -1613 -3357 -1603
rect -2858 -1610 -2857 -1600
rect -2855 -1610 -2853 -1600
rect -2849 -1610 -2847 -1600
rect -2845 -1610 -2844 -1600
rect -2229 -1601 -2227 -1591
rect -2225 -1601 -2215 -1591
rect -2904 -1620 -2902 -1610
rect -2900 -1620 -2890 -1610
rect -4136 -1663 -4134 -1653
rect -4132 -1663 -4122 -1653
rect -3663 -1658 -3662 -1638
rect -3660 -1658 -3652 -1638
rect -3650 -1658 -3649 -1638
rect -2810 -1613 -2808 -1603
rect -2806 -1613 -2796 -1603
rect -2135 -1594 -2133 -1584
rect -2131 -1594 -2121 -1584
rect -3614 -1655 -3612 -1645
rect -3610 -1655 -3600 -1645
rect -3817 -1678 -3815 -1668
rect -3813 -1678 -3803 -1668
rect -3769 -1678 -3768 -1668
rect -3766 -1678 -3764 -1668
rect -3760 -1678 -3758 -1668
rect -3756 -1678 -3755 -1668
rect -3721 -1681 -3719 -1671
rect -3717 -1681 -3707 -1671
rect -3311 -1656 -3310 -1636
rect -3308 -1656 -3300 -1636
rect -3298 -1656 -3297 -1636
rect -3262 -1653 -3260 -1643
rect -3258 -1653 -3248 -1643
rect -3465 -1676 -3463 -1666
rect -3461 -1676 -3451 -1666
rect -3417 -1676 -3416 -1666
rect -3414 -1676 -3412 -1666
rect -3408 -1676 -3406 -1666
rect -3404 -1676 -3403 -1666
rect -3369 -1679 -3367 -1669
rect -3365 -1679 -3355 -1669
rect -2750 -1656 -2749 -1636
rect -2747 -1656 -2739 -1636
rect -2737 -1656 -2736 -1636
rect -2075 -1637 -2074 -1617
rect -2072 -1637 -2064 -1617
rect -2062 -1637 -2061 -1617
rect -2026 -1634 -2024 -1624
rect -2022 -1634 -2012 -1624
rect -2701 -1653 -2699 -1643
rect -2697 -1653 -2687 -1643
rect -2904 -1676 -2902 -1666
rect -2900 -1676 -2890 -1666
rect -2856 -1676 -2855 -1666
rect -2853 -1676 -2851 -1666
rect -2847 -1676 -2845 -1666
rect -2843 -1676 -2842 -1666
rect -2808 -1679 -2806 -1669
rect -2804 -1679 -2794 -1669
rect -2229 -1657 -2227 -1647
rect -2225 -1657 -2215 -1647
rect -2181 -1657 -2180 -1647
rect -2178 -1657 -2176 -1647
rect -2172 -1657 -2170 -1647
rect -2168 -1657 -2167 -1647
rect -2133 -1660 -2131 -1650
rect -2129 -1660 -2119 -1650
rect -2194 -1736 -2193 -1726
rect -2191 -1736 -2189 -1726
rect -2185 -1736 -2183 -1726
rect -2181 -1736 -2180 -1726
rect -2146 -1739 -2144 -1729
rect -2142 -1739 -2132 -1729
rect -3414 -1767 -3413 -1757
rect -3411 -1767 -3409 -1757
rect -3405 -1767 -3403 -1757
rect -3401 -1767 -3400 -1757
rect -3801 -1787 -3800 -1777
rect -3798 -1787 -3796 -1777
rect -3792 -1787 -3790 -1777
rect -3788 -1787 -3787 -1777
rect -3753 -1790 -3751 -1780
rect -3749 -1790 -3739 -1780
rect -3366 -1770 -3364 -1760
rect -3362 -1770 -3352 -1760
rect -2864 -1766 -2863 -1756
rect -2861 -1766 -2859 -1756
rect -2855 -1766 -2853 -1756
rect -2851 -1766 -2850 -1756
rect -2816 -1769 -2814 -1759
rect -2812 -1769 -2802 -1759
rect -4247 -1841 -4246 -1821
rect -4244 -1841 -4238 -1821
rect -4236 -1841 -4235 -1821
rect -4195 -1841 -4194 -1831
rect -4192 -1841 -4191 -1831
rect -4161 -1834 -4160 -1824
rect -4158 -1834 -4157 -1824
rect -2948 -1844 -2947 -1824
rect -2945 -1844 -2939 -1824
rect -2937 -1844 -2936 -1824
rect -2896 -1844 -2895 -1834
rect -2893 -1844 -2892 -1834
rect -2862 -1837 -2861 -1827
rect -2859 -1837 -2858 -1827
rect -4117 -1854 -4115 -1844
rect -4113 -1854 -4103 -1844
rect -2710 -1840 -2709 -1820
rect -2707 -1840 -2701 -1820
rect -2699 -1840 -2698 -1820
rect -2658 -1840 -2657 -1830
rect -2655 -1840 -2654 -1830
rect -2624 -1833 -2623 -1823
rect -2621 -1833 -2620 -1823
rect -2261 -1829 -2260 -1809
rect -2258 -1829 -2252 -1809
rect -2250 -1829 -2249 -1809
rect -2209 -1829 -2208 -1819
rect -2206 -1829 -2205 -1819
rect -2175 -1822 -2174 -1812
rect -2172 -1822 -2171 -1812
rect -1944 -1822 -1943 -1802
rect -1941 -1822 -1935 -1802
rect -1933 -1822 -1932 -1802
rect -1892 -1822 -1891 -1812
rect -1889 -1822 -1888 -1812
rect -1858 -1815 -1857 -1805
rect -1855 -1815 -1854 -1805
rect -2818 -1857 -2816 -1847
rect -2814 -1857 -2804 -1847
rect -2580 -1853 -2578 -1843
rect -2576 -1853 -2566 -1843
rect -2131 -1842 -2129 -1832
rect -2127 -1842 -2117 -1832
rect -1814 -1835 -1812 -1825
rect -1810 -1835 -1800 -1825
rect -3623 -2002 -3622 -1982
rect -3620 -2002 -3614 -1982
rect -3612 -2002 -3611 -1982
rect -3571 -2002 -3570 -1992
rect -3568 -2002 -3567 -1992
rect -3537 -1995 -3536 -1985
rect -3534 -1995 -3533 -1985
rect -3324 -1993 -3323 -1973
rect -3321 -1993 -3315 -1973
rect -3313 -1993 -3312 -1973
rect -3272 -1993 -3271 -1983
rect -3269 -1993 -3268 -1983
rect -3238 -1986 -3237 -1976
rect -3235 -1986 -3234 -1976
rect -3493 -2015 -3491 -2005
rect -3489 -2015 -3479 -2005
rect -3194 -2006 -3192 -1996
rect -3190 -2006 -3180 -1996
<< ndcontact >>
rect -3291 -574 -3287 -569
rect -3275 -574 -3271 -569
rect -3851 -615 -3847 -610
rect -3835 -615 -3831 -610
rect -3247 -585 -3243 -575
rect -3224 -585 -3220 -575
rect -3205 -585 -3201 -575
rect -3189 -585 -3185 -575
rect -2292 -565 -2288 -560
rect -2276 -565 -2272 -560
rect -1662 -544 -1658 -539
rect -1646 -544 -1642 -539
rect -2248 -576 -2244 -566
rect -2225 -576 -2221 -566
rect -2206 -576 -2202 -566
rect -2190 -576 -2186 -566
rect -1618 -555 -1614 -545
rect -1595 -555 -1591 -545
rect -1576 -555 -1572 -545
rect -1560 -555 -1556 -545
rect -1532 -553 -1528 -548
rect -1514 -553 -1510 -548
rect -2162 -574 -2158 -569
rect -2144 -574 -2140 -569
rect -3161 -583 -3157 -578
rect -3143 -583 -3139 -578
rect -3807 -626 -3803 -616
rect -3784 -626 -3780 -616
rect -3765 -626 -3761 -616
rect -3749 -626 -3745 -616
rect -3721 -624 -3717 -619
rect -3703 -624 -3699 -619
rect -1931 -762 -1927 -757
rect -1913 -762 -1909 -757
rect -1885 -761 -1881 -751
rect -1867 -761 -1863 -751
rect -1837 -755 -1833 -750
rect -1819 -755 -1815 -750
rect -2553 -780 -2549 -775
rect -2535 -780 -2531 -775
rect -2507 -779 -2503 -769
rect -2489 -779 -2485 -769
rect -2459 -773 -2455 -768
rect -2441 -773 -2437 -768
rect -3274 -806 -3270 -801
rect -3256 -806 -3252 -801
rect -3228 -805 -3224 -795
rect -3210 -805 -3206 -795
rect -3180 -799 -3176 -794
rect -3162 -799 -3158 -794
rect -3274 -862 -3270 -857
rect -3256 -862 -3252 -857
rect -3071 -839 -3067 -834
rect -3053 -839 -3049 -834
rect -2553 -836 -2549 -831
rect -2535 -836 -2531 -831
rect -2350 -813 -2346 -808
rect -2332 -813 -2328 -808
rect -2399 -821 -2395 -816
rect -2391 -821 -2385 -816
rect -2381 -821 -2377 -816
rect -1931 -818 -1927 -813
rect -1913 -818 -1909 -813
rect -1728 -795 -1724 -790
rect -1710 -795 -1706 -790
rect -1777 -803 -1773 -798
rect -1769 -803 -1763 -798
rect -1759 -803 -1755 -798
rect -1883 -827 -1879 -817
rect -1865 -827 -1861 -817
rect -1835 -821 -1831 -816
rect -1817 -821 -1813 -816
rect -3120 -847 -3116 -842
rect -3112 -847 -3106 -842
rect -3102 -847 -3098 -842
rect -2505 -845 -2501 -835
rect -2487 -845 -2483 -835
rect -2457 -839 -2453 -834
rect -2439 -839 -2435 -834
rect -3226 -871 -3222 -861
rect -3208 -871 -3204 -861
rect -3178 -865 -3174 -860
rect -3160 -865 -3156 -860
rect -3819 -1052 -3815 -1047
rect -3801 -1052 -3797 -1047
rect -3773 -1051 -3769 -1041
rect -3755 -1051 -3751 -1041
rect -3725 -1045 -3721 -1040
rect -3707 -1045 -3703 -1040
rect -3819 -1108 -3815 -1103
rect -3801 -1108 -3797 -1103
rect -3616 -1085 -3612 -1080
rect -3598 -1085 -3594 -1080
rect -3665 -1093 -3661 -1088
rect -3657 -1093 -3651 -1088
rect -3647 -1093 -3643 -1088
rect -3771 -1117 -3767 -1107
rect -3753 -1117 -3749 -1107
rect -3723 -1111 -3719 -1106
rect -3705 -1111 -3701 -1106
rect -2433 -1157 -2429 -1147
rect -2415 -1157 -2411 -1147
rect -2385 -1151 -2381 -1146
rect -2367 -1151 -2363 -1146
rect -2245 -1204 -2241 -1199
rect -2227 -1204 -2223 -1199
rect -2294 -1212 -2290 -1207
rect -2286 -1212 -2280 -1207
rect -2276 -1212 -2272 -1207
rect -2434 -1280 -2430 -1270
rect -2416 -1280 -2412 -1270
rect -2386 -1274 -2382 -1269
rect -2368 -1274 -2364 -1269
rect -2918 -1313 -2914 -1303
rect -2900 -1313 -2896 -1303
rect -2870 -1307 -2866 -1302
rect -2852 -1307 -2848 -1302
rect -1884 -1315 -1880 -1310
rect -1866 -1315 -1862 -1310
rect -2069 -1324 -2065 -1319
rect -2051 -1324 -2047 -1319
rect -1933 -1323 -1929 -1318
rect -1925 -1323 -1919 -1318
rect -1915 -1323 -1911 -1318
rect -1824 -1319 -1820 -1314
rect -1808 -1319 -1804 -1314
rect -4304 -1363 -4300 -1358
rect -4288 -1363 -4284 -1358
rect -2118 -1332 -2114 -1327
rect -2110 -1332 -2104 -1327
rect -2100 -1332 -2096 -1327
rect -1780 -1330 -1776 -1320
rect -1757 -1330 -1753 -1320
rect -1738 -1330 -1734 -1320
rect -1722 -1330 -1718 -1320
rect -1694 -1328 -1690 -1323
rect -1676 -1328 -1672 -1323
rect -2737 -1349 -2733 -1344
rect -2719 -1349 -2715 -1344
rect -4260 -1374 -4256 -1364
rect -4237 -1374 -4233 -1364
rect -4218 -1374 -4214 -1364
rect -4202 -1374 -4198 -1364
rect -2786 -1357 -2782 -1352
rect -2778 -1357 -2772 -1352
rect -2768 -1357 -2764 -1352
rect -4174 -1372 -4170 -1367
rect -4156 -1372 -4152 -1367
rect -2621 -1388 -2617 -1383
rect -2603 -1388 -2599 -1383
rect -2670 -1396 -2666 -1391
rect -2662 -1396 -2656 -1391
rect -2652 -1396 -2648 -1391
rect -2429 -1403 -2425 -1393
rect -2411 -1403 -2407 -1393
rect -2381 -1397 -2377 -1392
rect -2363 -1397 -2359 -1392
rect -2919 -1419 -2915 -1409
rect -2901 -1419 -2897 -1409
rect -2871 -1413 -2867 -1408
rect -2853 -1413 -2849 -1408
rect -3490 -1430 -3486 -1420
rect -3472 -1430 -3468 -1420
rect -3442 -1424 -3438 -1419
rect -3424 -1424 -3420 -1419
rect -2733 -1451 -2729 -1446
rect -2715 -1451 -2711 -1446
rect -2246 -1448 -2242 -1443
rect -2228 -1448 -2224 -1443
rect -2782 -1459 -2778 -1454
rect -2774 -1459 -2768 -1454
rect -2764 -1459 -2760 -1454
rect -2295 -1456 -2291 -1451
rect -2287 -1456 -2281 -1451
rect -2277 -1456 -2273 -1451
rect -3200 -1482 -3196 -1477
rect -3182 -1482 -3178 -1477
rect -3315 -1492 -3311 -1487
rect -3297 -1492 -3293 -1487
rect -3249 -1490 -3245 -1485
rect -3241 -1490 -3235 -1485
rect -3231 -1490 -3227 -1485
rect -3364 -1500 -3360 -1495
rect -3356 -1500 -3350 -1495
rect -3346 -1500 -3342 -1495
rect -3824 -1548 -3820 -1538
rect -3806 -1548 -3802 -1538
rect -3776 -1542 -3772 -1537
rect -3758 -1542 -3754 -1537
rect -2915 -1516 -2911 -1506
rect -2897 -1516 -2893 -1506
rect -2867 -1510 -2863 -1505
rect -2849 -1510 -2845 -1505
rect -3671 -1540 -3667 -1535
rect -3653 -1540 -3649 -1535
rect -3485 -1539 -3481 -1529
rect -3467 -1539 -3463 -1529
rect -3437 -1533 -3433 -1528
rect -3419 -1533 -3415 -1528
rect -2430 -1531 -2426 -1521
rect -2412 -1531 -2408 -1521
rect -2382 -1525 -2378 -1520
rect -2364 -1525 -2360 -1520
rect -3720 -1548 -3716 -1543
rect -3712 -1548 -3706 -1543
rect -3702 -1548 -3698 -1543
rect -3821 -1642 -3817 -1637
rect -3803 -1642 -3799 -1637
rect -3775 -1641 -3771 -1631
rect -3757 -1641 -3753 -1631
rect -3727 -1635 -3723 -1630
rect -3709 -1635 -3705 -1630
rect -4270 -1674 -4266 -1669
rect -4254 -1674 -4250 -1669
rect -3469 -1640 -3465 -1635
rect -3451 -1640 -3447 -1635
rect -3423 -1639 -3419 -1629
rect -3405 -1639 -3401 -1629
rect -3375 -1633 -3371 -1628
rect -3357 -1633 -3353 -1628
rect -2233 -1621 -2229 -1616
rect -2215 -1621 -2211 -1616
rect -2187 -1620 -2183 -1610
rect -2169 -1620 -2165 -1610
rect -2139 -1614 -2135 -1609
rect -2121 -1614 -2117 -1609
rect -4226 -1685 -4222 -1675
rect -4203 -1685 -4199 -1675
rect -4184 -1685 -4180 -1675
rect -4168 -1685 -4164 -1675
rect -4140 -1683 -4136 -1678
rect -4122 -1683 -4118 -1678
rect -3821 -1698 -3817 -1693
rect -3803 -1698 -3799 -1693
rect -2908 -1640 -2904 -1635
rect -2890 -1640 -2886 -1635
rect -2862 -1639 -2858 -1629
rect -2844 -1639 -2840 -1629
rect -2814 -1633 -2810 -1628
rect -2796 -1633 -2792 -1628
rect -3618 -1675 -3614 -1670
rect -3600 -1675 -3596 -1670
rect -3667 -1683 -3663 -1678
rect -3659 -1683 -3653 -1678
rect -3649 -1683 -3645 -1678
rect -3469 -1696 -3465 -1691
rect -3451 -1696 -3447 -1691
rect -3266 -1673 -3262 -1668
rect -3248 -1673 -3244 -1668
rect -3315 -1681 -3311 -1676
rect -3307 -1681 -3301 -1676
rect -3297 -1681 -3293 -1676
rect -3773 -1707 -3769 -1697
rect -3755 -1707 -3751 -1697
rect -3725 -1701 -3721 -1696
rect -3707 -1701 -3703 -1696
rect -3421 -1705 -3417 -1695
rect -3403 -1705 -3399 -1695
rect -3373 -1699 -3369 -1694
rect -3355 -1699 -3351 -1694
rect -2908 -1696 -2904 -1691
rect -2890 -1696 -2886 -1691
rect -2705 -1673 -2701 -1668
rect -2687 -1673 -2683 -1668
rect -2754 -1681 -2750 -1676
rect -2746 -1681 -2740 -1676
rect -2736 -1681 -2732 -1676
rect -2233 -1677 -2229 -1672
rect -2215 -1677 -2211 -1672
rect -2030 -1654 -2026 -1649
rect -2012 -1654 -2008 -1649
rect -2079 -1662 -2075 -1657
rect -2071 -1662 -2065 -1657
rect -2061 -1662 -2057 -1657
rect -2185 -1686 -2181 -1676
rect -2167 -1686 -2163 -1676
rect -2137 -1680 -2133 -1675
rect -2119 -1680 -2115 -1675
rect -2860 -1705 -2856 -1695
rect -2842 -1705 -2838 -1695
rect -2812 -1699 -2808 -1694
rect -2794 -1699 -2790 -1694
rect -2198 -1765 -2194 -1755
rect -2180 -1765 -2176 -1755
rect -2150 -1759 -2146 -1754
rect -2132 -1759 -2128 -1754
rect -3418 -1796 -3414 -1786
rect -3400 -1796 -3396 -1786
rect -3370 -1790 -3366 -1785
rect -3352 -1790 -3348 -1785
rect -2868 -1795 -2864 -1785
rect -2850 -1795 -2846 -1785
rect -2820 -1789 -2816 -1784
rect -2802 -1789 -2798 -1784
rect -3805 -1816 -3801 -1806
rect -3787 -1816 -3783 -1806
rect -3757 -1810 -3753 -1805
rect -3739 -1810 -3735 -1805
rect -4251 -1865 -4247 -1860
rect -4235 -1865 -4231 -1860
rect -4207 -1876 -4203 -1866
rect -4184 -1876 -4180 -1866
rect -4165 -1876 -4161 -1866
rect -4149 -1876 -4145 -1866
rect -2952 -1868 -2948 -1863
rect -2936 -1868 -2932 -1863
rect -4121 -1874 -4117 -1869
rect -4103 -1874 -4099 -1869
rect -2908 -1879 -2904 -1869
rect -2885 -1879 -2881 -1869
rect -2866 -1879 -2862 -1869
rect -2850 -1879 -2846 -1869
rect -2714 -1864 -2710 -1859
rect -2698 -1864 -2694 -1859
rect -2265 -1853 -2261 -1848
rect -2249 -1853 -2245 -1848
rect -2822 -1877 -2818 -1872
rect -2804 -1877 -2800 -1872
rect -2670 -1875 -2666 -1865
rect -2647 -1875 -2643 -1865
rect -2628 -1875 -2624 -1865
rect -2612 -1875 -2608 -1865
rect -2221 -1864 -2217 -1854
rect -2198 -1864 -2194 -1854
rect -2179 -1864 -2175 -1854
rect -2163 -1864 -2159 -1854
rect -1948 -1846 -1944 -1841
rect -1932 -1846 -1928 -1841
rect -1904 -1857 -1900 -1847
rect -1881 -1857 -1877 -1847
rect -1862 -1857 -1858 -1847
rect -1846 -1857 -1842 -1847
rect -1818 -1855 -1814 -1850
rect -1800 -1855 -1796 -1850
rect -2135 -1862 -2131 -1857
rect -2117 -1862 -2113 -1857
rect -2584 -1873 -2580 -1868
rect -2566 -1873 -2562 -1868
rect -3627 -2026 -3623 -2021
rect -3611 -2026 -3607 -2021
rect -3583 -2037 -3579 -2027
rect -3560 -2037 -3556 -2027
rect -3541 -2037 -3537 -2027
rect -3525 -2037 -3521 -2027
rect -3328 -2017 -3324 -2012
rect -3312 -2017 -3308 -2012
rect -3284 -2028 -3280 -2018
rect -3261 -2028 -3257 -2018
rect -3242 -2028 -3238 -2018
rect -3226 -2028 -3222 -2018
rect -3198 -2026 -3194 -2021
rect -3180 -2026 -3176 -2021
rect -3497 -2035 -3493 -2030
rect -3479 -2035 -3475 -2030
<< pdcontact >>
rect -3291 -550 -3287 -530
rect -3275 -550 -3271 -530
rect -3239 -550 -3235 -540
rect -3231 -550 -3227 -540
rect -3205 -543 -3201 -533
rect -3197 -543 -3193 -533
rect -2292 -541 -2288 -521
rect -2276 -541 -2272 -521
rect -1662 -520 -1658 -500
rect -1646 -520 -1642 -500
rect -1610 -520 -1606 -510
rect -1602 -520 -1598 -510
rect -1576 -513 -1572 -503
rect -1568 -513 -1564 -503
rect -2240 -541 -2236 -531
rect -2232 -541 -2228 -531
rect -2206 -534 -2202 -524
rect -2198 -534 -2194 -524
rect -3851 -591 -3847 -571
rect -3835 -591 -3831 -571
rect -3799 -591 -3795 -581
rect -3791 -591 -3787 -581
rect -3765 -584 -3761 -574
rect -3757 -584 -3753 -574
rect -3161 -563 -3157 -553
rect -3143 -563 -3139 -553
rect -2162 -554 -2158 -544
rect -2144 -554 -2140 -544
rect -1532 -533 -1528 -523
rect -1514 -533 -1510 -523
rect -3721 -604 -3717 -594
rect -3703 -604 -3699 -594
rect -1885 -732 -1881 -722
rect -1876 -732 -1872 -722
rect -1867 -732 -1863 -722
rect -2507 -750 -2503 -740
rect -2498 -750 -2494 -740
rect -2489 -750 -2485 -740
rect -1931 -742 -1927 -732
rect -1913 -742 -1909 -732
rect -2553 -760 -2549 -750
rect -2535 -760 -2531 -750
rect -3228 -776 -3224 -766
rect -3219 -776 -3215 -766
rect -3210 -776 -3206 -766
rect -3274 -786 -3270 -776
rect -3256 -786 -3252 -776
rect -3180 -779 -3176 -769
rect -3162 -779 -3158 -769
rect -2459 -753 -2455 -743
rect -2441 -753 -2437 -743
rect -1837 -735 -1833 -725
rect -1819 -735 -1815 -725
rect -2399 -796 -2395 -776
rect -2381 -796 -2377 -776
rect -1777 -778 -1773 -758
rect -1759 -778 -1755 -758
rect -1728 -775 -1724 -765
rect -1710 -775 -1706 -765
rect -2350 -793 -2346 -783
rect -2332 -793 -2328 -783
rect -3120 -822 -3116 -802
rect -3102 -822 -3098 -802
rect -3071 -819 -3067 -809
rect -3053 -819 -3049 -809
rect -2553 -816 -2549 -806
rect -2535 -816 -2531 -806
rect -2505 -816 -2501 -806
rect -2496 -816 -2492 -806
rect -2487 -816 -2483 -806
rect -3274 -842 -3270 -832
rect -3256 -842 -3252 -832
rect -3226 -842 -3222 -832
rect -3217 -842 -3213 -832
rect -3208 -842 -3204 -832
rect -3178 -845 -3174 -835
rect -3160 -845 -3156 -835
rect -2457 -819 -2453 -809
rect -2439 -819 -2435 -809
rect -1931 -798 -1927 -788
rect -1913 -798 -1909 -788
rect -1883 -798 -1879 -788
rect -1874 -798 -1870 -788
rect -1865 -798 -1861 -788
rect -1835 -801 -1831 -791
rect -1817 -801 -1813 -791
rect -3773 -1022 -3769 -1012
rect -3764 -1022 -3760 -1012
rect -3755 -1022 -3751 -1012
rect -3819 -1032 -3815 -1022
rect -3801 -1032 -3797 -1022
rect -3725 -1025 -3721 -1015
rect -3707 -1025 -3703 -1015
rect -3665 -1068 -3661 -1048
rect -3647 -1068 -3643 -1048
rect -3616 -1065 -3612 -1055
rect -3598 -1065 -3594 -1055
rect -3819 -1088 -3815 -1078
rect -3801 -1088 -3797 -1078
rect -3771 -1088 -3767 -1078
rect -3762 -1088 -3758 -1078
rect -3753 -1088 -3749 -1078
rect -3723 -1091 -3719 -1081
rect -3705 -1091 -3701 -1081
rect -2433 -1128 -2429 -1118
rect -2424 -1128 -2420 -1118
rect -2415 -1128 -2411 -1118
rect -2385 -1131 -2381 -1121
rect -2367 -1131 -2363 -1121
rect -2294 -1187 -2290 -1167
rect -2276 -1187 -2272 -1167
rect -2245 -1184 -2241 -1174
rect -2227 -1184 -2223 -1174
rect -2434 -1251 -2430 -1241
rect -2425 -1251 -2421 -1241
rect -2416 -1251 -2412 -1241
rect -2386 -1254 -2382 -1244
rect -2368 -1254 -2364 -1244
rect -2918 -1284 -2914 -1274
rect -2909 -1284 -2905 -1274
rect -2900 -1284 -2896 -1274
rect -2870 -1287 -2866 -1277
rect -2852 -1287 -2848 -1277
rect -2118 -1307 -2114 -1287
rect -2100 -1307 -2096 -1287
rect -2069 -1304 -2065 -1294
rect -2051 -1304 -2047 -1294
rect -1933 -1298 -1929 -1278
rect -1915 -1298 -1911 -1278
rect -1884 -1295 -1880 -1285
rect -1866 -1295 -1862 -1285
rect -1824 -1295 -1820 -1275
rect -1808 -1295 -1804 -1275
rect -1772 -1295 -1768 -1285
rect -1764 -1295 -1760 -1285
rect -1738 -1288 -1734 -1278
rect -1730 -1288 -1726 -1278
rect -4304 -1339 -4300 -1319
rect -4288 -1339 -4284 -1319
rect -4252 -1339 -4248 -1329
rect -4244 -1339 -4240 -1329
rect -4218 -1332 -4214 -1322
rect -4210 -1332 -4206 -1322
rect -2786 -1332 -2782 -1312
rect -2768 -1332 -2764 -1312
rect -2737 -1329 -2733 -1319
rect -2719 -1329 -2715 -1319
rect -1694 -1308 -1690 -1298
rect -1676 -1308 -1672 -1298
rect -4174 -1352 -4170 -1342
rect -4156 -1352 -4152 -1342
rect -2670 -1371 -2666 -1351
rect -2652 -1371 -2648 -1351
rect -2621 -1368 -2617 -1358
rect -2603 -1368 -2599 -1358
rect -2919 -1390 -2915 -1380
rect -2910 -1390 -2906 -1380
rect -2901 -1390 -2897 -1380
rect -3490 -1401 -3486 -1391
rect -3481 -1401 -3477 -1391
rect -3472 -1401 -3468 -1391
rect -3442 -1404 -3438 -1394
rect -3424 -1404 -3420 -1394
rect -2871 -1393 -2867 -1383
rect -2853 -1393 -2849 -1383
rect -2429 -1374 -2425 -1364
rect -2420 -1374 -2416 -1364
rect -2411 -1374 -2407 -1364
rect -2381 -1377 -2377 -1367
rect -2363 -1377 -2359 -1367
rect -2782 -1434 -2778 -1414
rect -2764 -1434 -2760 -1414
rect -2733 -1431 -2729 -1421
rect -2715 -1431 -2711 -1421
rect -2295 -1431 -2291 -1411
rect -2277 -1431 -2273 -1411
rect -2246 -1428 -2242 -1418
rect -2228 -1428 -2224 -1418
rect -3364 -1475 -3360 -1455
rect -3346 -1475 -3342 -1455
rect -3315 -1472 -3311 -1462
rect -3297 -1472 -3293 -1462
rect -3249 -1465 -3245 -1445
rect -3231 -1465 -3227 -1445
rect -3200 -1462 -3196 -1452
rect -3182 -1462 -3178 -1452
rect -2915 -1487 -2911 -1477
rect -2906 -1487 -2902 -1477
rect -2897 -1487 -2893 -1477
rect -3824 -1519 -3820 -1509
rect -3815 -1519 -3811 -1509
rect -3806 -1519 -3802 -1509
rect -3776 -1522 -3772 -1512
rect -3758 -1522 -3754 -1512
rect -3720 -1523 -3716 -1503
rect -3702 -1523 -3698 -1503
rect -3485 -1510 -3481 -1500
rect -3476 -1510 -3472 -1500
rect -3467 -1510 -3463 -1500
rect -3671 -1520 -3667 -1510
rect -3653 -1520 -3649 -1510
rect -3437 -1513 -3433 -1503
rect -3419 -1513 -3415 -1503
rect -2867 -1490 -2863 -1480
rect -2849 -1490 -2845 -1480
rect -2430 -1502 -2426 -1492
rect -2421 -1502 -2417 -1492
rect -2412 -1502 -2408 -1492
rect -2382 -1505 -2378 -1495
rect -2364 -1505 -2360 -1495
rect -2187 -1591 -2183 -1581
rect -2178 -1591 -2174 -1581
rect -2169 -1591 -2165 -1581
rect -3775 -1612 -3771 -1602
rect -3766 -1612 -3762 -1602
rect -3757 -1612 -3753 -1602
rect -3821 -1622 -3817 -1612
rect -3803 -1622 -3799 -1612
rect -4270 -1650 -4266 -1630
rect -4254 -1650 -4250 -1630
rect -4218 -1650 -4214 -1640
rect -4210 -1650 -4206 -1640
rect -4184 -1643 -4180 -1633
rect -4176 -1643 -4172 -1633
rect -3727 -1615 -3723 -1605
rect -3709 -1615 -3705 -1605
rect -3423 -1610 -3419 -1600
rect -3414 -1610 -3410 -1600
rect -3405 -1610 -3401 -1600
rect -3469 -1620 -3465 -1610
rect -3451 -1620 -3447 -1610
rect -3375 -1613 -3371 -1603
rect -3357 -1613 -3353 -1603
rect -2862 -1610 -2858 -1600
rect -2853 -1610 -2849 -1600
rect -2844 -1610 -2840 -1600
rect -2233 -1601 -2229 -1591
rect -2215 -1601 -2211 -1591
rect -2908 -1620 -2904 -1610
rect -2890 -1620 -2886 -1610
rect -4140 -1663 -4136 -1653
rect -4122 -1663 -4118 -1653
rect -3667 -1658 -3663 -1638
rect -3649 -1658 -3645 -1638
rect -2814 -1613 -2810 -1603
rect -2796 -1613 -2792 -1603
rect -2139 -1594 -2135 -1584
rect -2121 -1594 -2117 -1584
rect -3618 -1655 -3614 -1645
rect -3600 -1655 -3596 -1645
rect -3821 -1678 -3817 -1668
rect -3803 -1678 -3799 -1668
rect -3773 -1678 -3769 -1668
rect -3764 -1678 -3760 -1668
rect -3755 -1678 -3751 -1668
rect -3725 -1681 -3721 -1671
rect -3707 -1681 -3703 -1671
rect -3315 -1656 -3311 -1636
rect -3297 -1656 -3293 -1636
rect -3266 -1653 -3262 -1643
rect -3248 -1653 -3244 -1643
rect -3469 -1676 -3465 -1666
rect -3451 -1676 -3447 -1666
rect -3421 -1676 -3417 -1666
rect -3412 -1676 -3408 -1666
rect -3403 -1676 -3399 -1666
rect -3373 -1679 -3369 -1669
rect -3355 -1679 -3351 -1669
rect -2754 -1656 -2750 -1636
rect -2736 -1656 -2732 -1636
rect -2079 -1637 -2075 -1617
rect -2061 -1637 -2057 -1617
rect -2030 -1634 -2026 -1624
rect -2012 -1634 -2008 -1624
rect -2705 -1653 -2701 -1643
rect -2687 -1653 -2683 -1643
rect -2908 -1676 -2904 -1666
rect -2890 -1676 -2886 -1666
rect -2860 -1676 -2856 -1666
rect -2851 -1676 -2847 -1666
rect -2842 -1676 -2838 -1666
rect -2812 -1679 -2808 -1669
rect -2794 -1679 -2790 -1669
rect -2233 -1657 -2229 -1647
rect -2215 -1657 -2211 -1647
rect -2185 -1657 -2181 -1647
rect -2176 -1657 -2172 -1647
rect -2167 -1657 -2163 -1647
rect -2137 -1660 -2133 -1650
rect -2119 -1660 -2115 -1650
rect -2198 -1736 -2194 -1726
rect -2189 -1736 -2185 -1726
rect -2180 -1736 -2176 -1726
rect -2150 -1739 -2146 -1729
rect -2132 -1739 -2128 -1729
rect -3418 -1767 -3414 -1757
rect -3409 -1767 -3405 -1757
rect -3400 -1767 -3396 -1757
rect -3805 -1787 -3801 -1777
rect -3796 -1787 -3792 -1777
rect -3787 -1787 -3783 -1777
rect -3757 -1790 -3753 -1780
rect -3739 -1790 -3735 -1780
rect -3370 -1770 -3366 -1760
rect -3352 -1770 -3348 -1760
rect -2868 -1766 -2864 -1756
rect -2859 -1766 -2855 -1756
rect -2850 -1766 -2846 -1756
rect -2820 -1769 -2816 -1759
rect -2802 -1769 -2798 -1759
rect -4251 -1841 -4247 -1821
rect -4235 -1841 -4231 -1821
rect -4199 -1841 -4195 -1831
rect -4191 -1841 -4187 -1831
rect -4165 -1834 -4161 -1824
rect -4157 -1834 -4153 -1824
rect -2952 -1844 -2948 -1824
rect -2936 -1844 -2932 -1824
rect -2900 -1844 -2896 -1834
rect -2892 -1844 -2888 -1834
rect -2866 -1837 -2862 -1827
rect -2858 -1837 -2854 -1827
rect -4121 -1854 -4117 -1844
rect -4103 -1854 -4099 -1844
rect -2714 -1840 -2710 -1820
rect -2698 -1840 -2694 -1820
rect -2662 -1840 -2658 -1830
rect -2654 -1840 -2650 -1830
rect -2628 -1833 -2624 -1823
rect -2620 -1833 -2616 -1823
rect -2265 -1829 -2261 -1809
rect -2249 -1829 -2245 -1809
rect -2213 -1829 -2209 -1819
rect -2205 -1829 -2201 -1819
rect -2179 -1822 -2175 -1812
rect -2171 -1822 -2167 -1812
rect -1948 -1822 -1944 -1802
rect -1932 -1822 -1928 -1802
rect -1896 -1822 -1892 -1812
rect -1888 -1822 -1884 -1812
rect -1862 -1815 -1858 -1805
rect -1854 -1815 -1850 -1805
rect -2822 -1857 -2818 -1847
rect -2804 -1857 -2800 -1847
rect -2584 -1853 -2580 -1843
rect -2566 -1853 -2562 -1843
rect -2135 -1842 -2131 -1832
rect -2117 -1842 -2113 -1832
rect -1818 -1835 -1814 -1825
rect -1800 -1835 -1796 -1825
rect -3627 -2002 -3623 -1982
rect -3611 -2002 -3607 -1982
rect -3575 -2002 -3571 -1992
rect -3567 -2002 -3563 -1992
rect -3541 -1995 -3537 -1985
rect -3533 -1995 -3529 -1985
rect -3328 -1993 -3324 -1973
rect -3312 -1993 -3308 -1973
rect -3276 -1993 -3272 -1983
rect -3268 -1993 -3264 -1983
rect -3242 -1986 -3238 -1976
rect -3234 -1986 -3230 -1976
rect -3497 -2015 -3493 -2005
rect -3479 -2015 -3475 -2005
rect -3198 -2006 -3194 -1996
rect -3180 -2006 -3176 -1996
<< polysilicon >>
rect -1657 -500 -1655 -497
rect -1649 -500 -1647 -497
rect -2287 -521 -2285 -518
rect -2279 -521 -2277 -518
rect -3286 -530 -3284 -527
rect -3278 -530 -3276 -527
rect -3234 -540 -3232 -532
rect -3200 -533 -3198 -528
rect -2235 -531 -2233 -523
rect -2201 -524 -2199 -519
rect -1605 -510 -1603 -502
rect -1571 -503 -1569 -498
rect -3846 -571 -3844 -568
rect -3838 -571 -3836 -568
rect -3286 -569 -3284 -550
rect -3278 -559 -3276 -550
rect -3278 -563 -3267 -559
rect -3794 -581 -3792 -573
rect -3760 -574 -3758 -569
rect -3242 -572 -3240 -567
rect -3286 -577 -3284 -574
rect -3234 -572 -3232 -550
rect -3200 -575 -3198 -543
rect -3155 -553 -3153 -550
rect -2287 -560 -2285 -541
rect -2279 -550 -2277 -541
rect -2279 -554 -2268 -550
rect -3192 -571 -3178 -567
rect -3192 -575 -3190 -571
rect -3846 -610 -3844 -591
rect -3838 -600 -3836 -591
rect -3838 -604 -3827 -600
rect -3802 -613 -3800 -608
rect -3846 -618 -3844 -615
rect -3794 -613 -3792 -591
rect -3760 -616 -3758 -584
rect -3155 -578 -3153 -563
rect -2243 -563 -2241 -558
rect -2287 -568 -2285 -565
rect -2235 -563 -2233 -541
rect -2201 -566 -2199 -534
rect -1657 -539 -1655 -520
rect -1649 -529 -1647 -520
rect -1649 -533 -1638 -529
rect -2156 -544 -2154 -541
rect -1613 -542 -1611 -537
rect -1657 -547 -1655 -544
rect -1605 -542 -1603 -520
rect -1571 -545 -1569 -513
rect -1526 -523 -1524 -520
rect -1563 -541 -1549 -537
rect -1563 -545 -1561 -541
rect -2193 -562 -2179 -558
rect -2193 -566 -2191 -562
rect -2156 -569 -2154 -554
rect -1526 -548 -1524 -533
rect -1613 -558 -1611 -555
rect -1605 -558 -1603 -555
rect -1571 -560 -1569 -555
rect -1563 -560 -1561 -555
rect -1526 -556 -1524 -553
rect -2243 -579 -2241 -576
rect -2235 -579 -2233 -576
rect -2201 -581 -2199 -576
rect -2193 -581 -2191 -576
rect -2156 -577 -2154 -574
rect -3242 -588 -3240 -585
rect -3234 -588 -3232 -585
rect -3200 -590 -3198 -585
rect -3192 -590 -3190 -585
rect -3155 -586 -3153 -583
rect -3715 -594 -3713 -591
rect -3752 -612 -3738 -608
rect -3752 -616 -3750 -612
rect -3715 -619 -3713 -604
rect -3802 -629 -3800 -626
rect -3794 -629 -3792 -626
rect -3760 -631 -3758 -626
rect -3752 -631 -3750 -626
rect -3715 -627 -3713 -624
rect -1880 -722 -1878 -719
rect -1870 -722 -1868 -719
rect -1925 -732 -1923 -729
rect -1831 -725 -1829 -722
rect -2502 -740 -2500 -737
rect -2492 -740 -2490 -737
rect -2547 -750 -2545 -747
rect -2453 -743 -2451 -740
rect -3223 -766 -3221 -763
rect -3213 -766 -3211 -763
rect -3268 -776 -3266 -773
rect -3174 -769 -3172 -766
rect -3268 -801 -3266 -786
rect -3223 -795 -3221 -776
rect -3213 -795 -3211 -776
rect -2547 -775 -2545 -760
rect -2502 -769 -2500 -750
rect -2492 -769 -2490 -750
rect -2453 -768 -2451 -753
rect -1925 -757 -1923 -742
rect -1880 -751 -1878 -732
rect -1870 -751 -1868 -732
rect -1831 -750 -1829 -735
rect -1831 -758 -1829 -755
rect -1772 -758 -1770 -755
rect -1762 -758 -1760 -755
rect -1925 -765 -1923 -762
rect -1880 -764 -1878 -761
rect -1870 -764 -1868 -761
rect -3174 -794 -3172 -779
rect -2453 -776 -2451 -773
rect -2394 -776 -2392 -773
rect -2384 -776 -2382 -773
rect -2547 -783 -2545 -780
rect -2502 -782 -2500 -779
rect -2492 -782 -2490 -779
rect -1722 -765 -1720 -762
rect -2344 -783 -2342 -780
rect -1925 -788 -1923 -785
rect -1878 -788 -1876 -785
rect -1868 -788 -1866 -785
rect -3174 -802 -3172 -799
rect -3115 -802 -3113 -799
rect -3105 -802 -3103 -799
rect -3268 -809 -3266 -806
rect -3223 -808 -3221 -805
rect -3213 -808 -3211 -805
rect -2547 -806 -2545 -803
rect -2500 -806 -2498 -803
rect -2490 -806 -2488 -803
rect -3065 -809 -3063 -806
rect -2451 -809 -2449 -806
rect -3268 -832 -3266 -829
rect -3221 -832 -3219 -829
rect -3211 -832 -3209 -829
rect -3172 -835 -3170 -832
rect -3268 -857 -3266 -842
rect -3221 -861 -3219 -842
rect -3211 -861 -3209 -842
rect -3115 -842 -3113 -822
rect -3105 -842 -3103 -822
rect -3065 -834 -3063 -819
rect -2547 -831 -2545 -816
rect -2500 -835 -2498 -816
rect -2490 -835 -2488 -816
rect -2394 -816 -2392 -796
rect -2384 -816 -2382 -796
rect -2344 -808 -2342 -793
rect -1829 -791 -1827 -788
rect -1925 -813 -1923 -798
rect -2344 -816 -2342 -813
rect -2451 -834 -2449 -819
rect -1878 -817 -1876 -798
rect -1868 -817 -1866 -798
rect -1772 -798 -1770 -778
rect -1762 -798 -1760 -778
rect -1722 -790 -1720 -775
rect -1722 -798 -1720 -795
rect -1829 -816 -1827 -801
rect -1772 -806 -1770 -803
rect -1762 -806 -1760 -803
rect -1925 -821 -1923 -818
rect -2394 -824 -2392 -821
rect -2384 -824 -2382 -821
rect -1829 -824 -1827 -821
rect -1878 -830 -1876 -827
rect -1868 -830 -1866 -827
rect -2547 -839 -2545 -836
rect -3065 -842 -3063 -839
rect -3172 -860 -3170 -845
rect -2451 -842 -2449 -839
rect -3115 -850 -3113 -847
rect -3105 -850 -3103 -847
rect -2500 -848 -2498 -845
rect -2490 -848 -2488 -845
rect -3268 -865 -3266 -862
rect -3172 -868 -3170 -865
rect -3221 -874 -3219 -871
rect -3211 -874 -3209 -871
rect -3768 -1012 -3766 -1009
rect -3758 -1012 -3756 -1009
rect -3813 -1022 -3811 -1019
rect -3719 -1015 -3717 -1012
rect -3813 -1047 -3811 -1032
rect -3768 -1041 -3766 -1022
rect -3758 -1041 -3756 -1022
rect -3719 -1040 -3717 -1025
rect -3719 -1048 -3717 -1045
rect -3660 -1048 -3658 -1045
rect -3650 -1048 -3648 -1045
rect -3813 -1055 -3811 -1052
rect -3768 -1054 -3766 -1051
rect -3758 -1054 -3756 -1051
rect -3610 -1055 -3608 -1052
rect -3813 -1078 -3811 -1075
rect -3766 -1078 -3764 -1075
rect -3756 -1078 -3754 -1075
rect -3717 -1081 -3715 -1078
rect -3813 -1103 -3811 -1088
rect -3766 -1107 -3764 -1088
rect -3756 -1107 -3754 -1088
rect -3660 -1088 -3658 -1068
rect -3650 -1088 -3648 -1068
rect -3610 -1080 -3608 -1065
rect -3610 -1088 -3608 -1085
rect -3717 -1106 -3715 -1091
rect -3660 -1096 -3658 -1093
rect -3650 -1096 -3648 -1093
rect -3813 -1111 -3811 -1108
rect -3717 -1114 -3715 -1111
rect -3766 -1120 -3764 -1117
rect -3756 -1120 -3754 -1117
rect -2428 -1118 -2426 -1115
rect -2418 -1118 -2416 -1115
rect -2379 -1121 -2377 -1118
rect -2428 -1147 -2426 -1128
rect -2418 -1147 -2416 -1128
rect -2379 -1146 -2377 -1131
rect -2379 -1154 -2377 -1151
rect -2428 -1160 -2426 -1157
rect -2418 -1160 -2416 -1157
rect -2289 -1167 -2287 -1164
rect -2279 -1167 -2277 -1164
rect -2239 -1174 -2237 -1171
rect -2289 -1207 -2287 -1187
rect -2279 -1207 -2277 -1187
rect -2239 -1199 -2237 -1184
rect -2239 -1207 -2237 -1204
rect -2289 -1215 -2287 -1212
rect -2279 -1215 -2277 -1212
rect -2429 -1241 -2427 -1238
rect -2419 -1241 -2417 -1238
rect -2380 -1244 -2378 -1241
rect -2429 -1270 -2427 -1251
rect -2419 -1270 -2417 -1251
rect -2380 -1269 -2378 -1254
rect -2913 -1274 -2911 -1271
rect -2903 -1274 -2901 -1271
rect -2864 -1277 -2862 -1274
rect -2913 -1303 -2911 -1284
rect -2903 -1303 -2901 -1284
rect -2380 -1277 -2378 -1274
rect -1819 -1275 -1817 -1272
rect -1811 -1275 -1809 -1272
rect -1928 -1278 -1926 -1275
rect -1918 -1278 -1916 -1275
rect -2429 -1283 -2427 -1280
rect -2419 -1283 -2417 -1280
rect -2113 -1287 -2111 -1284
rect -2103 -1287 -2101 -1284
rect -2864 -1302 -2862 -1287
rect -2063 -1294 -2061 -1291
rect -1878 -1285 -1876 -1282
rect -1767 -1285 -1765 -1277
rect -1733 -1278 -1731 -1273
rect -2864 -1310 -2862 -1307
rect -2781 -1312 -2779 -1309
rect -2771 -1312 -2769 -1309
rect -2913 -1316 -2911 -1313
rect -2903 -1316 -2901 -1313
rect -4299 -1319 -4297 -1316
rect -4291 -1319 -4289 -1316
rect -4247 -1329 -4245 -1321
rect -4213 -1322 -4211 -1317
rect -2731 -1319 -2729 -1316
rect -2113 -1327 -2111 -1307
rect -2103 -1327 -2101 -1307
rect -2063 -1319 -2061 -1304
rect -1928 -1318 -1926 -1298
rect -1918 -1318 -1916 -1298
rect -1878 -1310 -1876 -1295
rect -1819 -1314 -1817 -1295
rect -1811 -1304 -1809 -1295
rect -1811 -1308 -1800 -1304
rect -1878 -1318 -1876 -1315
rect -1775 -1317 -1773 -1312
rect -1819 -1322 -1817 -1319
rect -1767 -1317 -1765 -1295
rect -1733 -1320 -1731 -1288
rect -1688 -1298 -1686 -1295
rect -1725 -1316 -1711 -1312
rect -1725 -1320 -1723 -1316
rect -2063 -1327 -2061 -1324
rect -1928 -1326 -1926 -1323
rect -1918 -1326 -1916 -1323
rect -4299 -1358 -4297 -1339
rect -4291 -1348 -4289 -1339
rect -4291 -1352 -4280 -1348
rect -4255 -1361 -4253 -1356
rect -4299 -1366 -4297 -1363
rect -4247 -1361 -4245 -1339
rect -4213 -1364 -4211 -1332
rect -4168 -1342 -4166 -1339
rect -2781 -1352 -2779 -1332
rect -2771 -1352 -2769 -1332
rect -2731 -1344 -2729 -1329
rect -1688 -1323 -1686 -1308
rect -2113 -1335 -2111 -1332
rect -2103 -1335 -2101 -1332
rect -1775 -1333 -1773 -1330
rect -1767 -1333 -1765 -1330
rect -1733 -1335 -1731 -1330
rect -1725 -1335 -1723 -1330
rect -1688 -1331 -1686 -1328
rect -2731 -1352 -2729 -1349
rect -2665 -1351 -2663 -1348
rect -2655 -1351 -2653 -1348
rect -4205 -1360 -4191 -1356
rect -4205 -1364 -4203 -1360
rect -4168 -1367 -4166 -1352
rect -2781 -1360 -2779 -1357
rect -2771 -1360 -2769 -1357
rect -2615 -1358 -2613 -1355
rect -2424 -1364 -2422 -1361
rect -2414 -1364 -2412 -1361
rect -4255 -1377 -4253 -1374
rect -4247 -1377 -4245 -1374
rect -4213 -1379 -4211 -1374
rect -4205 -1379 -4203 -1374
rect -4168 -1375 -4166 -1372
rect -2914 -1380 -2912 -1377
rect -2904 -1380 -2902 -1377
rect -3485 -1391 -3483 -1388
rect -3475 -1391 -3473 -1388
rect -2865 -1383 -2863 -1380
rect -3436 -1394 -3434 -1391
rect -3485 -1420 -3483 -1401
rect -3475 -1420 -3473 -1401
rect -3436 -1419 -3434 -1404
rect -2914 -1409 -2912 -1390
rect -2904 -1409 -2902 -1390
rect -2665 -1391 -2663 -1371
rect -2655 -1391 -2653 -1371
rect -2615 -1383 -2613 -1368
rect -2375 -1367 -2373 -1364
rect -2615 -1391 -2613 -1388
rect -2865 -1408 -2863 -1393
rect -2424 -1393 -2422 -1374
rect -2414 -1393 -2412 -1374
rect -2375 -1392 -2373 -1377
rect -2665 -1399 -2663 -1396
rect -2655 -1399 -2653 -1396
rect -2375 -1400 -2373 -1397
rect -2424 -1406 -2422 -1403
rect -2414 -1406 -2412 -1403
rect -2290 -1411 -2288 -1408
rect -2280 -1411 -2278 -1408
rect -2865 -1416 -2863 -1413
rect -2777 -1414 -2775 -1411
rect -2767 -1414 -2765 -1411
rect -2914 -1422 -2912 -1419
rect -2904 -1422 -2902 -1419
rect -3436 -1427 -3434 -1424
rect -3485 -1433 -3483 -1430
rect -3475 -1433 -3473 -1430
rect -2727 -1421 -2725 -1418
rect -2240 -1418 -2238 -1415
rect -3244 -1445 -3242 -1442
rect -3234 -1445 -3232 -1442
rect -3359 -1455 -3357 -1452
rect -3349 -1455 -3347 -1452
rect -3309 -1462 -3307 -1459
rect -3194 -1452 -3192 -1449
rect -2777 -1454 -2775 -1434
rect -2767 -1454 -2765 -1434
rect -2727 -1446 -2725 -1431
rect -2290 -1451 -2288 -1431
rect -2280 -1451 -2278 -1431
rect -2240 -1443 -2238 -1428
rect -2240 -1451 -2238 -1448
rect -2727 -1454 -2725 -1451
rect -2290 -1459 -2288 -1456
rect -2280 -1459 -2278 -1456
rect -2777 -1462 -2775 -1459
rect -2767 -1462 -2765 -1459
rect -3359 -1495 -3357 -1475
rect -3349 -1495 -3347 -1475
rect -3309 -1487 -3307 -1472
rect -3244 -1485 -3242 -1465
rect -3234 -1485 -3232 -1465
rect -3194 -1477 -3192 -1462
rect -2910 -1477 -2908 -1474
rect -2900 -1477 -2898 -1474
rect -3194 -1485 -3192 -1482
rect -2861 -1480 -2859 -1477
rect -3309 -1495 -3307 -1492
rect -3244 -1493 -3242 -1490
rect -3234 -1493 -3232 -1490
rect -3480 -1500 -3478 -1497
rect -3470 -1500 -3468 -1497
rect -3715 -1503 -3713 -1500
rect -3705 -1503 -3703 -1500
rect -3819 -1509 -3817 -1506
rect -3809 -1509 -3807 -1506
rect -3770 -1512 -3768 -1509
rect -3819 -1538 -3817 -1519
rect -3809 -1538 -3807 -1519
rect -3770 -1537 -3768 -1522
rect -3665 -1510 -3663 -1507
rect -3431 -1503 -3429 -1500
rect -3359 -1503 -3357 -1500
rect -3349 -1503 -3347 -1500
rect -3770 -1545 -3768 -1542
rect -3715 -1543 -3713 -1523
rect -3705 -1543 -3703 -1523
rect -3665 -1535 -3663 -1520
rect -3480 -1529 -3478 -1510
rect -3470 -1529 -3468 -1510
rect -2910 -1506 -2908 -1487
rect -2900 -1506 -2898 -1487
rect -2861 -1505 -2859 -1490
rect -2425 -1492 -2423 -1489
rect -2415 -1492 -2413 -1489
rect -2376 -1495 -2374 -1492
rect -3431 -1528 -3429 -1513
rect -2861 -1513 -2859 -1510
rect -2910 -1519 -2908 -1516
rect -2900 -1519 -2898 -1516
rect -2425 -1521 -2423 -1502
rect -2415 -1521 -2413 -1502
rect -2376 -1520 -2374 -1505
rect -2376 -1528 -2374 -1525
rect -3431 -1536 -3429 -1533
rect -2425 -1534 -2423 -1531
rect -2415 -1534 -2413 -1531
rect -3665 -1543 -3663 -1540
rect -3480 -1542 -3478 -1539
rect -3470 -1542 -3468 -1539
rect -3819 -1551 -3817 -1548
rect -3809 -1551 -3807 -1548
rect -3715 -1551 -3713 -1548
rect -3705 -1551 -3703 -1548
rect -2182 -1581 -2180 -1578
rect -2172 -1581 -2170 -1578
rect -2227 -1591 -2225 -1588
rect -2133 -1584 -2131 -1581
rect -3770 -1602 -3768 -1599
rect -3760 -1602 -3758 -1599
rect -3418 -1600 -3416 -1597
rect -3408 -1600 -3406 -1597
rect -2857 -1600 -2855 -1597
rect -2847 -1600 -2845 -1597
rect -3815 -1612 -3813 -1609
rect -3721 -1605 -3719 -1602
rect -4265 -1630 -4263 -1627
rect -4257 -1630 -4255 -1627
rect -4213 -1640 -4211 -1632
rect -4179 -1633 -4177 -1628
rect -3815 -1637 -3813 -1622
rect -3770 -1631 -3768 -1612
rect -3760 -1631 -3758 -1612
rect -3463 -1610 -3461 -1607
rect -3369 -1603 -3367 -1600
rect -3721 -1630 -3719 -1615
rect -3463 -1635 -3461 -1620
rect -3418 -1629 -3416 -1610
rect -3408 -1629 -3406 -1610
rect -2902 -1610 -2900 -1607
rect -2808 -1603 -2806 -1600
rect -3369 -1628 -3367 -1613
rect -3721 -1638 -3719 -1635
rect -3662 -1638 -3660 -1635
rect -3652 -1638 -3650 -1635
rect -4265 -1669 -4263 -1650
rect -4257 -1659 -4255 -1650
rect -4257 -1663 -4246 -1659
rect -4221 -1672 -4219 -1667
rect -4265 -1677 -4263 -1674
rect -4213 -1672 -4211 -1650
rect -4179 -1675 -4177 -1643
rect -3815 -1645 -3813 -1642
rect -3770 -1644 -3768 -1641
rect -3760 -1644 -3758 -1641
rect -4134 -1653 -4132 -1650
rect -3369 -1636 -3367 -1633
rect -3310 -1636 -3308 -1633
rect -3300 -1636 -3298 -1633
rect -2902 -1635 -2900 -1620
rect -2857 -1629 -2855 -1610
rect -2847 -1629 -2845 -1610
rect -2808 -1628 -2806 -1613
rect -2227 -1616 -2225 -1601
rect -2182 -1610 -2180 -1591
rect -2172 -1610 -2170 -1591
rect -2133 -1609 -2131 -1594
rect -2133 -1617 -2131 -1614
rect -2074 -1617 -2072 -1614
rect -2064 -1617 -2062 -1614
rect -2227 -1624 -2225 -1621
rect -2182 -1623 -2180 -1620
rect -2172 -1623 -2170 -1620
rect -3612 -1645 -3610 -1642
rect -3463 -1643 -3461 -1640
rect -3418 -1642 -3416 -1639
rect -3408 -1642 -3406 -1639
rect -4171 -1671 -4157 -1667
rect -4171 -1675 -4169 -1671
rect -4134 -1678 -4132 -1663
rect -3815 -1668 -3813 -1665
rect -3768 -1668 -3766 -1665
rect -3758 -1668 -3756 -1665
rect -3719 -1671 -3717 -1668
rect -4221 -1688 -4219 -1685
rect -4213 -1688 -4211 -1685
rect -4179 -1690 -4177 -1685
rect -4171 -1690 -4169 -1685
rect -4134 -1686 -4132 -1683
rect -3815 -1693 -3813 -1678
rect -3768 -1697 -3766 -1678
rect -3758 -1697 -3756 -1678
rect -3662 -1678 -3660 -1658
rect -3652 -1678 -3650 -1658
rect -3612 -1670 -3610 -1655
rect -2808 -1636 -2806 -1633
rect -2749 -1636 -2747 -1633
rect -2739 -1636 -2737 -1633
rect -3260 -1643 -3258 -1640
rect -2902 -1643 -2900 -1640
rect -2857 -1642 -2855 -1639
rect -2847 -1642 -2845 -1639
rect -3463 -1666 -3461 -1663
rect -3416 -1666 -3414 -1663
rect -3406 -1666 -3404 -1663
rect -3612 -1678 -3610 -1675
rect -3367 -1669 -3365 -1666
rect -3719 -1696 -3717 -1681
rect -3662 -1686 -3660 -1683
rect -3652 -1686 -3650 -1683
rect -3463 -1691 -3461 -1676
rect -3416 -1695 -3414 -1676
rect -3406 -1695 -3404 -1676
rect -3310 -1676 -3308 -1656
rect -3300 -1676 -3298 -1656
rect -3260 -1668 -3258 -1653
rect -2024 -1624 -2022 -1621
rect -2699 -1643 -2697 -1640
rect -2227 -1647 -2225 -1644
rect -2180 -1647 -2178 -1644
rect -2170 -1647 -2168 -1644
rect -2902 -1666 -2900 -1663
rect -2855 -1666 -2853 -1663
rect -2845 -1666 -2843 -1663
rect -3260 -1676 -3258 -1673
rect -2806 -1669 -2804 -1666
rect -3367 -1694 -3365 -1679
rect -3310 -1684 -3308 -1681
rect -3300 -1684 -3298 -1681
rect -2902 -1691 -2900 -1676
rect -3815 -1701 -3813 -1698
rect -3463 -1699 -3461 -1696
rect -3719 -1704 -3717 -1701
rect -2855 -1695 -2853 -1676
rect -2845 -1695 -2843 -1676
rect -2749 -1676 -2747 -1656
rect -2739 -1676 -2737 -1656
rect -2699 -1668 -2697 -1653
rect -2131 -1650 -2129 -1647
rect -2227 -1672 -2225 -1657
rect -2699 -1676 -2697 -1673
rect -2806 -1694 -2804 -1679
rect -2180 -1676 -2178 -1657
rect -2170 -1676 -2168 -1657
rect -2074 -1657 -2072 -1637
rect -2064 -1657 -2062 -1637
rect -2024 -1649 -2022 -1634
rect -2024 -1657 -2022 -1654
rect -2131 -1675 -2129 -1660
rect -2074 -1665 -2072 -1662
rect -2064 -1665 -2062 -1662
rect -2227 -1680 -2225 -1677
rect -2749 -1684 -2747 -1681
rect -2739 -1684 -2737 -1681
rect -2131 -1683 -2129 -1680
rect -2180 -1689 -2178 -1686
rect -2170 -1689 -2168 -1686
rect -2902 -1699 -2900 -1696
rect -3367 -1702 -3365 -1699
rect -2806 -1702 -2804 -1699
rect -3768 -1710 -3766 -1707
rect -3758 -1710 -3756 -1707
rect -3416 -1708 -3414 -1705
rect -3406 -1708 -3404 -1705
rect -2855 -1708 -2853 -1705
rect -2845 -1708 -2843 -1705
rect -2193 -1726 -2191 -1723
rect -2183 -1726 -2181 -1723
rect -2144 -1729 -2142 -1726
rect -3413 -1757 -3411 -1754
rect -3403 -1757 -3401 -1754
rect -2863 -1756 -2861 -1753
rect -2853 -1756 -2851 -1753
rect -2193 -1755 -2191 -1736
rect -2183 -1755 -2181 -1736
rect -2144 -1754 -2142 -1739
rect -3364 -1760 -3362 -1757
rect -3800 -1777 -3798 -1774
rect -3790 -1777 -3788 -1774
rect -3751 -1780 -3749 -1777
rect -3800 -1806 -3798 -1787
rect -3790 -1806 -3788 -1787
rect -3413 -1786 -3411 -1767
rect -3403 -1786 -3401 -1767
rect -2814 -1759 -2812 -1756
rect -3364 -1785 -3362 -1770
rect -2863 -1785 -2861 -1766
rect -2853 -1785 -2851 -1766
rect -2144 -1762 -2142 -1759
rect -2193 -1768 -2191 -1765
rect -2183 -1768 -2181 -1765
rect -2814 -1784 -2812 -1769
rect -3751 -1805 -3749 -1790
rect -3364 -1793 -3362 -1790
rect -2814 -1792 -2812 -1789
rect -3413 -1799 -3411 -1796
rect -3403 -1799 -3401 -1796
rect -2863 -1798 -2861 -1795
rect -2853 -1798 -2851 -1795
rect -1943 -1802 -1941 -1799
rect -1935 -1802 -1933 -1799
rect -2260 -1809 -2258 -1806
rect -2252 -1809 -2250 -1806
rect -3751 -1813 -3749 -1810
rect -4246 -1821 -4244 -1818
rect -4238 -1821 -4236 -1818
rect -3800 -1819 -3798 -1816
rect -3790 -1819 -3788 -1816
rect -4194 -1831 -4192 -1823
rect -4160 -1824 -4158 -1819
rect -2709 -1820 -2707 -1817
rect -2701 -1820 -2699 -1817
rect -2947 -1824 -2945 -1821
rect -2939 -1824 -2937 -1821
rect -4246 -1860 -4244 -1841
rect -4238 -1850 -4236 -1841
rect -4238 -1854 -4227 -1850
rect -4202 -1863 -4200 -1858
rect -4246 -1868 -4244 -1865
rect -4194 -1863 -4192 -1841
rect -4160 -1866 -4158 -1834
rect -4115 -1844 -4113 -1841
rect -2895 -1834 -2893 -1826
rect -2861 -1827 -2859 -1822
rect -4152 -1862 -4138 -1858
rect -4152 -1866 -4150 -1862
rect -4115 -1869 -4113 -1854
rect -2947 -1863 -2945 -1844
rect -2939 -1853 -2937 -1844
rect -2939 -1857 -2928 -1853
rect -2903 -1866 -2901 -1861
rect -2947 -1871 -2945 -1868
rect -2895 -1866 -2893 -1844
rect -2861 -1869 -2859 -1837
rect -2657 -1830 -2655 -1822
rect -2623 -1823 -2621 -1818
rect -2208 -1819 -2206 -1811
rect -2174 -1812 -2172 -1807
rect -1891 -1812 -1889 -1804
rect -1857 -1805 -1855 -1800
rect -2816 -1847 -2814 -1844
rect -2853 -1865 -2839 -1861
rect -2853 -1869 -2851 -1865
rect -4202 -1879 -4200 -1876
rect -4194 -1879 -4192 -1876
rect -4160 -1881 -4158 -1876
rect -4152 -1881 -4150 -1876
rect -4115 -1877 -4113 -1874
rect -2816 -1872 -2814 -1857
rect -2709 -1859 -2707 -1840
rect -2701 -1849 -2699 -1840
rect -2701 -1853 -2690 -1849
rect -2665 -1862 -2663 -1857
rect -2709 -1867 -2707 -1864
rect -2657 -1862 -2655 -1840
rect -2623 -1865 -2621 -1833
rect -2578 -1843 -2576 -1840
rect -2260 -1848 -2258 -1829
rect -2252 -1838 -2250 -1829
rect -2252 -1842 -2241 -1838
rect -2216 -1851 -2214 -1846
rect -2615 -1861 -2601 -1857
rect -2615 -1865 -2613 -1861
rect -2578 -1868 -2576 -1853
rect -2260 -1856 -2258 -1853
rect -2208 -1851 -2206 -1829
rect -2174 -1854 -2172 -1822
rect -2129 -1832 -2127 -1829
rect -1943 -1841 -1941 -1822
rect -1935 -1831 -1933 -1822
rect -1935 -1835 -1924 -1831
rect -2166 -1850 -2152 -1846
rect -2166 -1854 -2164 -1850
rect -2129 -1857 -2127 -1842
rect -1899 -1844 -1897 -1839
rect -1943 -1849 -1941 -1846
rect -1891 -1844 -1889 -1822
rect -1857 -1847 -1855 -1815
rect -1812 -1825 -1810 -1822
rect -1849 -1843 -1835 -1839
rect -1849 -1847 -1847 -1843
rect -1812 -1850 -1810 -1835
rect -1899 -1860 -1897 -1857
rect -1891 -1860 -1889 -1857
rect -1857 -1862 -1855 -1857
rect -1849 -1862 -1847 -1857
rect -1812 -1858 -1810 -1855
rect -2216 -1867 -2214 -1864
rect -2208 -1867 -2206 -1864
rect -2174 -1869 -2172 -1864
rect -2166 -1869 -2164 -1864
rect -2129 -1865 -2127 -1862
rect -2903 -1882 -2901 -1879
rect -2895 -1882 -2893 -1879
rect -2861 -1884 -2859 -1879
rect -2853 -1884 -2851 -1879
rect -2816 -1880 -2814 -1877
rect -2665 -1878 -2663 -1875
rect -2657 -1878 -2655 -1875
rect -2623 -1880 -2621 -1875
rect -2615 -1880 -2613 -1875
rect -2578 -1876 -2576 -1873
rect -3323 -1973 -3321 -1970
rect -3315 -1973 -3313 -1970
rect -3622 -1982 -3620 -1979
rect -3614 -1982 -3612 -1979
rect -3570 -1992 -3568 -1984
rect -3536 -1985 -3534 -1980
rect -3271 -1983 -3269 -1975
rect -3237 -1976 -3235 -1971
rect -3622 -2021 -3620 -2002
rect -3614 -2011 -3612 -2002
rect -3614 -2015 -3603 -2011
rect -3578 -2024 -3576 -2019
rect -3622 -2029 -3620 -2026
rect -3570 -2024 -3568 -2002
rect -3536 -2027 -3534 -1995
rect -3491 -2005 -3489 -2002
rect -3323 -2012 -3321 -1993
rect -3315 -2002 -3313 -1993
rect -3315 -2006 -3304 -2002
rect -3528 -2023 -3514 -2019
rect -3528 -2027 -3526 -2023
rect -3491 -2030 -3489 -2015
rect -3279 -2015 -3277 -2010
rect -3323 -2020 -3321 -2017
rect -3271 -2015 -3269 -1993
rect -3237 -2018 -3235 -1986
rect -3192 -1996 -3190 -1993
rect -3229 -2014 -3215 -2010
rect -3229 -2018 -3227 -2014
rect -3192 -2021 -3190 -2006
rect -3279 -2031 -3277 -2028
rect -3271 -2031 -3269 -2028
rect -3237 -2033 -3235 -2028
rect -3229 -2033 -3227 -2028
rect -3192 -2029 -3190 -2026
rect -3578 -2040 -3576 -2037
rect -3570 -2040 -3568 -2037
rect -3536 -2042 -3534 -2037
rect -3528 -2042 -3526 -2037
rect -3491 -2038 -3489 -2035
<< polycontact >>
rect -1661 -532 -1657 -528
rect -3290 -562 -3286 -558
rect -3267 -563 -3263 -559
rect -3238 -563 -3234 -559
rect -3247 -572 -3242 -567
rect -3204 -572 -3200 -568
rect -2291 -553 -2287 -549
rect -2268 -554 -2264 -550
rect -2239 -554 -2235 -550
rect -3182 -567 -3178 -563
rect -3159 -575 -3155 -571
rect -3850 -603 -3846 -599
rect -3827 -604 -3823 -600
rect -3798 -604 -3794 -600
rect -3807 -613 -3802 -608
rect -3764 -613 -3760 -609
rect -2248 -563 -2243 -558
rect -2205 -563 -2201 -559
rect -1638 -533 -1634 -529
rect -1609 -533 -1605 -529
rect -1618 -542 -1613 -537
rect -1575 -542 -1571 -538
rect -1553 -537 -1549 -533
rect -1530 -545 -1526 -541
rect -2183 -558 -2179 -554
rect -2160 -566 -2156 -562
rect -3742 -608 -3738 -604
rect -3719 -616 -3715 -612
rect -3272 -798 -3268 -794
rect -3227 -787 -3223 -783
rect -2551 -772 -2547 -768
rect -2506 -761 -2502 -757
rect -2490 -761 -2486 -757
rect -2457 -765 -2453 -761
rect -1929 -754 -1925 -750
rect -1884 -743 -1880 -739
rect -1868 -743 -1864 -739
rect -1835 -747 -1831 -743
rect -3211 -787 -3207 -783
rect -3178 -791 -3174 -787
rect -2398 -807 -2394 -803
rect -3119 -833 -3115 -829
rect -3272 -854 -3268 -850
rect -3225 -853 -3221 -849
rect -3109 -833 -3105 -829
rect -3069 -831 -3065 -827
rect -2551 -828 -2547 -824
rect -2504 -827 -2500 -823
rect -2388 -807 -2384 -803
rect -2348 -805 -2344 -801
rect -1776 -789 -1772 -785
rect -1929 -810 -1925 -806
rect -1882 -809 -1878 -805
rect -2488 -827 -2484 -823
rect -2455 -831 -2451 -827
rect -1766 -789 -1762 -785
rect -1726 -787 -1722 -783
rect -1866 -809 -1862 -805
rect -1833 -813 -1829 -809
rect -3209 -853 -3205 -849
rect -3176 -857 -3172 -853
rect -3817 -1044 -3813 -1040
rect -3772 -1033 -3768 -1029
rect -3756 -1033 -3752 -1029
rect -3723 -1037 -3719 -1033
rect -3664 -1079 -3660 -1075
rect -3817 -1100 -3813 -1096
rect -3770 -1099 -3766 -1095
rect -3654 -1079 -3650 -1075
rect -3614 -1077 -3610 -1073
rect -3754 -1099 -3750 -1095
rect -3721 -1103 -3717 -1099
rect -2432 -1140 -2428 -1135
rect -2416 -1139 -2412 -1135
rect -2383 -1143 -2379 -1139
rect -2293 -1198 -2289 -1194
rect -2283 -1198 -2279 -1194
rect -2243 -1196 -2239 -1192
rect -2433 -1262 -2429 -1258
rect -2417 -1262 -2413 -1258
rect -2384 -1266 -2380 -1262
rect -2917 -1295 -2913 -1291
rect -2901 -1295 -2897 -1291
rect -2868 -1299 -2864 -1295
rect -2117 -1318 -2113 -1314
rect -2107 -1318 -2103 -1314
rect -2067 -1316 -2063 -1312
rect -1932 -1309 -1928 -1305
rect -1922 -1309 -1918 -1305
rect -1882 -1307 -1878 -1303
rect -1823 -1307 -1819 -1303
rect -1800 -1308 -1796 -1304
rect -1771 -1308 -1767 -1304
rect -1780 -1317 -1775 -1312
rect -1737 -1317 -1733 -1313
rect -1715 -1312 -1711 -1308
rect -1692 -1320 -1688 -1316
rect -4303 -1351 -4299 -1347
rect -4280 -1352 -4276 -1348
rect -4251 -1352 -4247 -1348
rect -4260 -1361 -4255 -1356
rect -4217 -1361 -4213 -1357
rect -2785 -1343 -2781 -1339
rect -2775 -1343 -2771 -1339
rect -2735 -1341 -2731 -1337
rect -4195 -1356 -4191 -1352
rect -4172 -1364 -4168 -1360
rect -2669 -1382 -2665 -1378
rect -3489 -1413 -3485 -1408
rect -2918 -1401 -2914 -1397
rect -3473 -1412 -3469 -1408
rect -3440 -1416 -3436 -1412
rect -2659 -1382 -2655 -1378
rect -2619 -1380 -2615 -1376
rect -2428 -1385 -2424 -1381
rect -2902 -1401 -2898 -1397
rect -2869 -1405 -2865 -1401
rect -2412 -1385 -2408 -1381
rect -2379 -1389 -2375 -1385
rect -2781 -1445 -2777 -1441
rect -2771 -1445 -2767 -1441
rect -2731 -1443 -2727 -1439
rect -2294 -1442 -2290 -1438
rect -2284 -1442 -2280 -1438
rect -2244 -1440 -2240 -1436
rect -3363 -1486 -3359 -1482
rect -3353 -1486 -3349 -1482
rect -3313 -1484 -3309 -1480
rect -3248 -1476 -3244 -1472
rect -3238 -1476 -3234 -1472
rect -3198 -1474 -3194 -1470
rect -2914 -1498 -2910 -1494
rect -3823 -1530 -3819 -1526
rect -3807 -1530 -3803 -1526
rect -3774 -1534 -3770 -1530
rect -3719 -1534 -3715 -1530
rect -3709 -1534 -3705 -1530
rect -3669 -1532 -3665 -1528
rect -3484 -1521 -3480 -1517
rect -2898 -1498 -2894 -1494
rect -2865 -1502 -2861 -1498
rect -3468 -1521 -3464 -1517
rect -3435 -1525 -3431 -1521
rect -2429 -1513 -2425 -1509
rect -2413 -1513 -2409 -1509
rect -2380 -1517 -2376 -1513
rect -3819 -1634 -3815 -1630
rect -3774 -1623 -3770 -1619
rect -3758 -1623 -3754 -1619
rect -3725 -1627 -3721 -1623
rect -3467 -1632 -3463 -1628
rect -3422 -1621 -3418 -1617
rect -3406 -1621 -3402 -1617
rect -3373 -1625 -3369 -1621
rect -4269 -1662 -4265 -1658
rect -4246 -1663 -4242 -1659
rect -4217 -1663 -4213 -1659
rect -4226 -1672 -4221 -1667
rect -4183 -1672 -4179 -1668
rect -2906 -1632 -2902 -1627
rect -2861 -1621 -2857 -1617
rect -2231 -1613 -2227 -1609
rect -2845 -1621 -2841 -1617
rect -2812 -1625 -2808 -1621
rect -2186 -1602 -2182 -1598
rect -2170 -1602 -2166 -1598
rect -2137 -1606 -2133 -1602
rect -4161 -1667 -4157 -1663
rect -4138 -1675 -4134 -1671
rect -3666 -1669 -3662 -1665
rect -3819 -1690 -3815 -1686
rect -3772 -1689 -3768 -1685
rect -3656 -1669 -3652 -1665
rect -3616 -1667 -3612 -1663
rect -3314 -1667 -3310 -1663
rect -3756 -1689 -3752 -1685
rect -3723 -1693 -3719 -1689
rect -3467 -1688 -3463 -1684
rect -3420 -1687 -3416 -1683
rect -3304 -1667 -3300 -1663
rect -3264 -1665 -3260 -1661
rect -2753 -1667 -2749 -1663
rect -3404 -1687 -3400 -1683
rect -3371 -1691 -3367 -1687
rect -2906 -1688 -2902 -1684
rect -2859 -1687 -2855 -1683
rect -2743 -1667 -2739 -1663
rect -2703 -1665 -2699 -1661
rect -2078 -1648 -2074 -1644
rect -2231 -1669 -2227 -1665
rect -2184 -1668 -2180 -1664
rect -2843 -1687 -2839 -1683
rect -2810 -1691 -2806 -1687
rect -2068 -1648 -2064 -1644
rect -2028 -1646 -2024 -1642
rect -2168 -1668 -2164 -1664
rect -2135 -1672 -2131 -1668
rect -2197 -1747 -2193 -1743
rect -2181 -1747 -2177 -1743
rect -2148 -1751 -2144 -1747
rect -3417 -1779 -3413 -1774
rect -3804 -1799 -3800 -1794
rect -3401 -1778 -3397 -1774
rect -3368 -1782 -3364 -1778
rect -2867 -1778 -2863 -1773
rect -2851 -1777 -2847 -1773
rect -2818 -1781 -2814 -1777
rect -3788 -1798 -3784 -1794
rect -3755 -1802 -3751 -1798
rect -4250 -1853 -4246 -1849
rect -4227 -1854 -4223 -1850
rect -4198 -1854 -4194 -1850
rect -4207 -1863 -4202 -1858
rect -4164 -1863 -4160 -1859
rect -4142 -1858 -4138 -1854
rect -4119 -1866 -4115 -1862
rect -2951 -1856 -2947 -1852
rect -2928 -1857 -2924 -1853
rect -2899 -1857 -2895 -1853
rect -2908 -1866 -2903 -1861
rect -2865 -1866 -2861 -1862
rect -2713 -1852 -2709 -1848
rect -2843 -1861 -2839 -1857
rect -2820 -1869 -2816 -1865
rect -2690 -1853 -2686 -1849
rect -2661 -1853 -2657 -1849
rect -2670 -1862 -2665 -1857
rect -2627 -1862 -2623 -1858
rect -2264 -1841 -2260 -1837
rect -2241 -1842 -2237 -1838
rect -2212 -1842 -2208 -1838
rect -2221 -1851 -2216 -1846
rect -2605 -1857 -2601 -1853
rect -2582 -1865 -2578 -1861
rect -2178 -1851 -2174 -1847
rect -1947 -1834 -1943 -1830
rect -1924 -1835 -1920 -1831
rect -1895 -1835 -1891 -1831
rect -2156 -1846 -2152 -1842
rect -2133 -1854 -2129 -1850
rect -1904 -1844 -1899 -1839
rect -1861 -1844 -1857 -1840
rect -1839 -1839 -1835 -1835
rect -1816 -1847 -1812 -1843
rect -3626 -2014 -3622 -2010
rect -3603 -2015 -3599 -2011
rect -3574 -2015 -3570 -2011
rect -3583 -2024 -3578 -2019
rect -3540 -2024 -3536 -2020
rect -3327 -2005 -3323 -2001
rect -3304 -2006 -3300 -2002
rect -3275 -2006 -3271 -2002
rect -3518 -2019 -3514 -2015
rect -3495 -2027 -3491 -2023
rect -3284 -2015 -3279 -2010
rect -3241 -2015 -3237 -2011
rect -3219 -2010 -3215 -2006
rect -3196 -2018 -3192 -2014
<< polynplus >>
rect -3242 -575 -3240 -572
rect -3234 -575 -3232 -572
rect -3802 -616 -3800 -613
rect -3794 -616 -3792 -613
rect -2243 -566 -2241 -563
rect -2235 -566 -2233 -563
rect -1613 -545 -1611 -542
rect -1605 -545 -1603 -542
rect -1775 -1320 -1773 -1317
rect -1767 -1320 -1765 -1317
rect -4255 -1364 -4253 -1361
rect -4247 -1364 -4245 -1361
rect -4221 -1675 -4219 -1672
rect -4213 -1675 -4211 -1672
rect -4202 -1866 -4200 -1863
rect -4194 -1866 -4192 -1863
rect -2903 -1869 -2901 -1866
rect -2895 -1869 -2893 -1866
rect -2665 -1865 -2663 -1862
rect -2657 -1865 -2655 -1862
rect -2216 -1854 -2214 -1851
rect -2208 -1854 -2206 -1851
rect -1899 -1847 -1897 -1844
rect -1891 -1847 -1889 -1844
rect -3578 -2027 -3576 -2024
rect -3570 -2027 -3568 -2024
rect -3279 -2018 -3277 -2015
rect -3271 -2018 -3269 -2015
<< metal1 >>
rect -1668 -496 -1636 -493
rect -1616 -496 -1592 -493
rect -1582 -496 -1558 -493
rect -1662 -500 -1658 -496
rect -2298 -517 -2266 -514
rect -2246 -517 -2222 -514
rect -2212 -517 -2188 -514
rect -2292 -521 -2288 -517
rect -3297 -526 -3265 -523
rect -3245 -526 -3221 -523
rect -3211 -526 -3187 -523
rect -3291 -530 -3287 -526
rect -3239 -540 -3235 -526
rect -3205 -533 -3201 -526
rect -2240 -531 -2236 -517
rect -2206 -524 -2202 -517
rect -1610 -510 -1606 -496
rect -1576 -503 -1572 -496
rect -3857 -567 -3825 -564
rect -3805 -567 -3781 -564
rect -3771 -567 -3747 -564
rect -3851 -571 -3847 -567
rect -3799 -581 -3795 -567
rect -3765 -574 -3761 -567
rect -3275 -569 -3271 -550
rect -3268 -569 -3247 -567
rect -3271 -572 -3247 -569
rect -3231 -568 -3227 -550
rect -3197 -561 -3193 -543
rect -3167 -547 -3133 -543
rect -3161 -553 -3157 -547
rect -3197 -565 -3185 -561
rect -2276 -560 -2272 -541
rect -2269 -560 -2248 -558
rect -3231 -572 -3204 -568
rect -3189 -571 -3185 -565
rect -3143 -571 -3139 -563
rect -2272 -563 -2248 -560
rect -2232 -559 -2228 -541
rect -2198 -552 -2194 -534
rect -2168 -538 -2134 -534
rect -2162 -544 -2158 -538
rect -1646 -539 -1642 -520
rect -1639 -539 -1618 -537
rect -1642 -542 -1618 -539
rect -1602 -538 -1598 -520
rect -1568 -531 -1564 -513
rect -1538 -517 -1504 -513
rect -1532 -523 -1528 -517
rect -1568 -535 -1556 -531
rect -1602 -542 -1575 -538
rect -1560 -541 -1556 -535
rect -1514 -541 -1510 -533
rect -1642 -544 -1634 -542
rect -2198 -556 -2186 -552
rect -1662 -549 -1658 -544
rect -1668 -552 -1636 -549
rect -2232 -563 -2205 -559
rect -2190 -562 -2186 -556
rect -2144 -562 -2140 -554
rect -1618 -561 -1614 -555
rect -1602 -561 -1598 -542
rect -1560 -545 -1530 -541
rect -1514 -545 -1504 -541
rect -2272 -565 -2264 -563
rect -2292 -570 -2288 -565
rect -3271 -574 -3263 -572
rect -3291 -579 -3287 -574
rect -3297 -582 -3265 -579
rect -3835 -610 -3831 -591
rect -3828 -610 -3807 -608
rect -3831 -613 -3807 -610
rect -3791 -609 -3787 -591
rect -3757 -602 -3753 -584
rect -3727 -588 -3693 -584
rect -3721 -594 -3717 -588
rect -3247 -591 -3243 -585
rect -3231 -591 -3227 -572
rect -3189 -575 -3159 -571
rect -3143 -575 -3133 -571
rect -2298 -573 -2266 -570
rect -3757 -606 -3745 -602
rect -3247 -595 -3227 -591
rect -3224 -598 -3220 -585
rect -3143 -578 -3139 -575
rect -2248 -582 -2244 -576
rect -2232 -582 -2228 -563
rect -2190 -566 -2160 -562
rect -2144 -566 -2134 -562
rect -1618 -565 -1598 -561
rect -3205 -596 -3201 -585
rect -3161 -589 -3157 -583
rect -2248 -586 -2228 -582
rect -2225 -589 -2221 -576
rect -2144 -569 -2140 -566
rect -1595 -568 -1591 -555
rect -1514 -548 -1510 -545
rect -1576 -566 -1572 -555
rect -1532 -559 -1528 -553
rect -1538 -562 -1504 -559
rect -1621 -573 -1587 -568
rect -1579 -571 -1555 -566
rect -2206 -587 -2202 -576
rect -2162 -580 -2158 -574
rect -2168 -583 -2134 -580
rect -3167 -592 -3133 -589
rect -2251 -594 -2217 -589
rect -2209 -592 -2185 -587
rect -3250 -603 -3216 -598
rect -3208 -601 -3184 -596
rect -3791 -613 -3764 -609
rect -3749 -612 -3745 -606
rect -3703 -611 -3699 -604
rect -3831 -615 -3823 -613
rect -3851 -620 -3847 -615
rect -3857 -623 -3825 -620
rect -3807 -632 -3803 -626
rect -3791 -632 -3787 -613
rect -3749 -616 -3719 -612
rect -3703 -616 -3678 -611
rect -3807 -636 -3787 -632
rect -3784 -639 -3780 -626
rect -3703 -619 -3699 -616
rect -3765 -637 -3761 -626
rect -3721 -630 -3717 -624
rect -3727 -633 -3693 -630
rect -3810 -644 -3776 -639
rect -3768 -642 -3744 -637
rect -1891 -717 -1857 -713
rect -1885 -722 -1881 -717
rect -1867 -722 -1863 -717
rect -1843 -719 -1809 -715
rect -1937 -726 -1903 -722
rect -2513 -735 -2479 -731
rect -1931 -732 -1927 -726
rect -1837 -725 -1833 -719
rect -2507 -740 -2503 -735
rect -2489 -740 -2485 -735
rect -2465 -737 -2431 -733
rect -2559 -744 -2525 -740
rect -2553 -750 -2549 -744
rect -2459 -743 -2455 -737
rect -3234 -761 -3200 -757
rect -2644 -759 -2574 -752
rect -3228 -766 -3224 -761
rect -3210 -766 -3206 -761
rect -3186 -763 -3152 -759
rect -3280 -770 -3246 -766
rect -3274 -776 -3270 -770
rect -3180 -769 -3176 -763
rect -3330 -783 -3295 -778
rect -3330 -806 -3325 -783
rect -3304 -794 -3301 -793
rect -3256 -794 -3252 -786
rect -3243 -787 -3227 -783
rect -3243 -794 -3239 -787
rect -3219 -790 -3215 -776
rect -3207 -787 -3203 -783
rect -3162 -787 -3158 -779
rect -3219 -791 -3206 -790
rect -3193 -791 -3178 -787
rect -3162 -791 -3142 -787
rect -3219 -794 -3189 -791
rect -3162 -794 -3158 -791
rect -3304 -798 -3272 -794
rect -3256 -798 -3239 -794
rect -3210 -795 -3189 -794
rect -3256 -801 -3252 -798
rect -4012 -811 -3325 -806
rect -3180 -805 -3176 -799
rect -4012 -1271 -4007 -811
rect -3274 -812 -3270 -806
rect -3228 -809 -3224 -805
rect -3186 -808 -3152 -805
rect -3234 -812 -3200 -809
rect -3280 -815 -3246 -812
rect -3280 -826 -3246 -822
rect -3274 -832 -3270 -826
rect -3232 -827 -3198 -823
rect -3226 -832 -3222 -827
rect -3208 -832 -3204 -827
rect -3184 -829 -3150 -825
rect -3147 -829 -3142 -791
rect -3126 -794 -3092 -790
rect -3120 -802 -3116 -794
rect -3077 -803 -3043 -799
rect -3071 -809 -3067 -803
rect -3178 -835 -3174 -829
rect -3147 -833 -3119 -829
rect -3102 -835 -3098 -822
rect -3053 -826 -3049 -819
rect -3089 -831 -3069 -827
rect -3053 -831 -3036 -826
rect -3089 -835 -3085 -831
rect -3053 -834 -3049 -831
rect -3256 -850 -3252 -842
rect -3242 -850 -3225 -849
rect -3288 -854 -3272 -850
rect -3256 -853 -3225 -850
rect -3256 -854 -3241 -853
rect -3256 -857 -3252 -854
rect -3217 -856 -3213 -842
rect -3102 -836 -3085 -835
rect -3112 -839 -3085 -836
rect -3112 -842 -3106 -839
rect -3205 -853 -3201 -849
rect -3160 -853 -3156 -845
rect -3071 -845 -3067 -839
rect -3217 -857 -3204 -856
rect -3191 -857 -3176 -853
rect -3160 -857 -3146 -853
rect -3120 -853 -3116 -847
rect -3102 -853 -3098 -847
rect -3077 -848 -3043 -845
rect -3126 -856 -3092 -853
rect -3217 -860 -3187 -857
rect -3160 -860 -3156 -857
rect -3208 -861 -3187 -860
rect -3274 -868 -3270 -862
rect -3280 -871 -3246 -868
rect -3178 -871 -3174 -865
rect -3226 -875 -3222 -871
rect -3184 -874 -3150 -871
rect -3232 -878 -3201 -875
rect -2644 -982 -2635 -759
rect -2583 -768 -2580 -767
rect -2535 -768 -2531 -760
rect -2522 -761 -2506 -757
rect -2522 -768 -2518 -761
rect -2498 -764 -2494 -750
rect -2486 -761 -2482 -757
rect -2441 -761 -2437 -753
rect -1961 -750 -1958 -749
rect -1913 -750 -1909 -742
rect -1900 -743 -1884 -739
rect -1900 -750 -1896 -743
rect -1876 -746 -1872 -732
rect -1864 -743 -1860 -739
rect -1819 -743 -1815 -735
rect -1876 -747 -1863 -746
rect -1850 -747 -1835 -743
rect -1819 -747 -1799 -743
rect -1876 -750 -1846 -747
rect -1819 -750 -1815 -747
rect -1961 -754 -1929 -750
rect -1913 -754 -1896 -750
rect -1867 -751 -1846 -750
rect -1913 -757 -1909 -754
rect -2498 -765 -2485 -764
rect -2472 -765 -2457 -761
rect -2441 -765 -2421 -761
rect -1837 -761 -1833 -755
rect -2498 -768 -2468 -765
rect -2441 -768 -2437 -765
rect -2583 -772 -2551 -768
rect -2535 -772 -2518 -768
rect -2489 -769 -2468 -768
rect -2535 -775 -2531 -772
rect -2459 -779 -2455 -773
rect -2553 -786 -2549 -780
rect -2507 -783 -2503 -779
rect -2465 -782 -2431 -779
rect -2513 -786 -2479 -783
rect -2559 -789 -2525 -786
rect -2559 -800 -2525 -796
rect -2553 -806 -2549 -800
rect -2511 -801 -2477 -797
rect -2505 -806 -2501 -801
rect -2487 -806 -2483 -801
rect -2463 -803 -2429 -799
rect -2426 -803 -2421 -765
rect -2405 -768 -2371 -764
rect -1931 -768 -1927 -762
rect -1885 -765 -1881 -761
rect -1843 -764 -1809 -761
rect -1891 -768 -1857 -765
rect -2399 -776 -2395 -768
rect -1937 -771 -1903 -768
rect -2356 -777 -2322 -773
rect -2350 -783 -2346 -777
rect -1937 -782 -1903 -778
rect -2457 -809 -2453 -803
rect -2426 -807 -2398 -803
rect -2381 -809 -2377 -796
rect -2332 -800 -2328 -793
rect -1931 -788 -1927 -782
rect -1889 -783 -1855 -779
rect -1883 -788 -1879 -783
rect -1865 -788 -1861 -783
rect -1841 -785 -1807 -781
rect -1804 -785 -1799 -747
rect -1783 -750 -1749 -746
rect -1777 -758 -1773 -750
rect -1734 -759 -1700 -755
rect -1728 -765 -1724 -759
rect -1835 -791 -1831 -785
rect -1804 -789 -1776 -785
rect -1759 -791 -1755 -778
rect -1710 -782 -1706 -775
rect -1746 -787 -1726 -783
rect -1710 -787 -1687 -782
rect -1746 -791 -1742 -787
rect -1710 -790 -1706 -787
rect -2368 -805 -2348 -801
rect -2332 -805 -2311 -800
rect -2368 -809 -2364 -805
rect -2332 -808 -2328 -805
rect -2535 -824 -2531 -816
rect -2521 -824 -2504 -823
rect -2567 -828 -2551 -824
rect -2535 -827 -2504 -824
rect -2535 -828 -2520 -827
rect -2535 -831 -2531 -828
rect -2496 -830 -2492 -816
rect -2381 -810 -2364 -809
rect -2391 -813 -2364 -810
rect -1913 -806 -1909 -798
rect -1899 -806 -1882 -805
rect -1945 -810 -1929 -806
rect -1913 -809 -1882 -806
rect -1913 -810 -1898 -809
rect -1913 -813 -1909 -810
rect -2391 -816 -2385 -813
rect -2484 -827 -2480 -823
rect -2439 -827 -2435 -819
rect -2350 -819 -2346 -813
rect -1874 -812 -1870 -798
rect -1759 -792 -1742 -791
rect -1769 -795 -1742 -792
rect -1769 -798 -1763 -795
rect -1728 -801 -1724 -795
rect -1862 -809 -1858 -805
rect -1777 -809 -1773 -803
rect -1759 -809 -1755 -803
rect -1734 -804 -1700 -801
rect -1874 -813 -1861 -812
rect -1848 -813 -1833 -809
rect -1783 -812 -1749 -809
rect -1874 -816 -1844 -813
rect -1865 -817 -1844 -816
rect -2496 -831 -2483 -830
rect -2470 -831 -2455 -827
rect -2439 -831 -2425 -827
rect -2399 -827 -2395 -821
rect -2381 -827 -2377 -821
rect -2356 -822 -2322 -819
rect -1931 -824 -1927 -818
rect -1937 -827 -1903 -824
rect -1835 -827 -1831 -821
rect -2405 -830 -2371 -827
rect -1883 -831 -1879 -827
rect -1841 -830 -1807 -827
rect -2496 -834 -2466 -831
rect -2439 -834 -2435 -831
rect -1889 -834 -1858 -831
rect -2487 -835 -2466 -834
rect -2553 -842 -2549 -836
rect -2559 -845 -2525 -842
rect -2457 -845 -2453 -839
rect -2505 -849 -2501 -845
rect -2463 -848 -2429 -845
rect -2511 -852 -2480 -849
rect -3012 -986 -2635 -982
rect -3155 -987 -2636 -986
rect -3155 -991 -3007 -987
rect -3779 -1007 -3745 -1003
rect -3773 -1012 -3769 -1007
rect -3755 -1012 -3751 -1007
rect -3731 -1009 -3697 -1005
rect -3825 -1016 -3791 -1012
rect -3819 -1022 -3815 -1016
rect -3725 -1015 -3721 -1009
rect -3936 -1271 -3931 -1032
rect -3849 -1040 -3846 -1039
rect -3801 -1040 -3797 -1032
rect -3788 -1033 -3772 -1029
rect -3788 -1040 -3784 -1033
rect -3764 -1036 -3760 -1022
rect -3752 -1033 -3748 -1029
rect -3707 -1033 -3703 -1025
rect -3764 -1037 -3751 -1036
rect -3738 -1037 -3723 -1033
rect -3707 -1037 -3687 -1033
rect -3764 -1040 -3734 -1037
rect -3707 -1040 -3703 -1037
rect -3849 -1044 -3817 -1040
rect -3801 -1044 -3784 -1040
rect -3755 -1041 -3734 -1040
rect -3801 -1047 -3797 -1044
rect -3725 -1051 -3721 -1045
rect -3819 -1058 -3815 -1052
rect -3773 -1055 -3769 -1051
rect -3731 -1054 -3697 -1051
rect -3779 -1058 -3745 -1055
rect -3825 -1061 -3791 -1058
rect -3825 -1072 -3791 -1068
rect -3819 -1078 -3815 -1072
rect -3777 -1073 -3743 -1069
rect -3771 -1078 -3767 -1073
rect -3753 -1078 -3749 -1073
rect -3729 -1075 -3695 -1071
rect -3692 -1075 -3687 -1037
rect -3671 -1040 -3637 -1036
rect -3665 -1048 -3661 -1040
rect -3622 -1049 -3588 -1045
rect -3616 -1055 -3612 -1049
rect -3723 -1081 -3719 -1075
rect -3692 -1079 -3664 -1075
rect -3647 -1081 -3643 -1068
rect -3598 -1072 -3594 -1065
rect -3634 -1077 -3614 -1073
rect -3598 -1077 -3552 -1072
rect -3634 -1081 -3630 -1077
rect -3598 -1080 -3594 -1077
rect -3801 -1096 -3797 -1088
rect -3787 -1096 -3770 -1095
rect -3833 -1100 -3817 -1096
rect -3801 -1099 -3770 -1096
rect -3801 -1100 -3786 -1099
rect -3801 -1103 -3797 -1100
rect -3762 -1102 -3758 -1088
rect -3647 -1082 -3630 -1081
rect -3657 -1085 -3630 -1082
rect -3657 -1088 -3651 -1085
rect -3750 -1099 -3746 -1095
rect -3705 -1099 -3701 -1091
rect -3616 -1091 -3612 -1085
rect -3762 -1103 -3749 -1102
rect -3736 -1103 -3721 -1099
rect -3705 -1103 -3691 -1099
rect -3665 -1099 -3661 -1093
rect -3647 -1099 -3643 -1093
rect -3622 -1094 -3588 -1091
rect -3671 -1102 -3637 -1099
rect -3762 -1106 -3732 -1103
rect -3705 -1106 -3701 -1103
rect -3753 -1107 -3732 -1106
rect -3819 -1114 -3815 -1108
rect -3825 -1117 -3791 -1114
rect -3723 -1117 -3719 -1111
rect -3771 -1121 -3767 -1117
rect -3729 -1120 -3695 -1117
rect -3777 -1124 -3746 -1121
rect -4310 -1315 -4278 -1312
rect -4258 -1315 -4234 -1312
rect -4224 -1315 -4200 -1312
rect -4304 -1319 -4300 -1315
rect -4252 -1329 -4248 -1315
rect -4218 -1322 -4214 -1315
rect -4288 -1358 -4284 -1339
rect -4281 -1358 -4260 -1356
rect -4284 -1361 -4260 -1358
rect -4244 -1357 -4240 -1339
rect -4210 -1350 -4206 -1332
rect -4180 -1336 -4146 -1332
rect -4174 -1342 -4170 -1336
rect -4210 -1354 -4198 -1350
rect -4244 -1361 -4217 -1357
rect -4202 -1360 -4198 -1354
rect -4156 -1359 -4152 -1352
rect -4284 -1363 -4276 -1361
rect -4304 -1368 -4300 -1363
rect -4310 -1371 -4278 -1368
rect -4260 -1380 -4256 -1374
rect -4244 -1380 -4240 -1361
rect -4202 -1364 -4172 -1360
rect -4156 -1364 -4131 -1359
rect -4260 -1384 -4240 -1380
rect -4237 -1387 -4233 -1374
rect -4156 -1367 -4152 -1364
rect -4218 -1385 -4214 -1374
rect -4174 -1378 -4170 -1372
rect -4180 -1381 -4146 -1378
rect -4263 -1392 -4229 -1387
rect -4221 -1390 -4197 -1385
rect -4276 -1626 -4244 -1623
rect -4224 -1626 -4200 -1623
rect -4190 -1626 -4166 -1623
rect -4270 -1630 -4266 -1626
rect -4218 -1640 -4214 -1626
rect -4184 -1633 -4180 -1626
rect -4254 -1669 -4250 -1650
rect -4247 -1669 -4226 -1667
rect -4250 -1672 -4226 -1669
rect -4210 -1668 -4206 -1650
rect -4176 -1661 -4172 -1643
rect -4146 -1647 -4112 -1643
rect -4140 -1653 -4136 -1647
rect -4176 -1665 -4164 -1661
rect -4210 -1672 -4183 -1668
rect -4168 -1671 -4164 -1665
rect -4122 -1670 -4118 -1663
rect -4250 -1674 -4242 -1672
rect -4270 -1679 -4266 -1674
rect -4276 -1682 -4244 -1679
rect -4226 -1691 -4222 -1685
rect -4210 -1691 -4206 -1672
rect -4168 -1675 -4138 -1671
rect -4122 -1675 -4095 -1670
rect -4226 -1695 -4206 -1691
rect -4203 -1698 -4199 -1685
rect -4122 -1678 -4118 -1675
rect -4184 -1696 -4180 -1685
rect -4140 -1689 -4136 -1683
rect -4146 -1692 -4112 -1689
rect -4229 -1703 -4195 -1698
rect -4187 -1701 -4163 -1696
rect -4257 -1817 -4225 -1814
rect -4205 -1817 -4181 -1814
rect -4171 -1817 -4147 -1814
rect -4251 -1821 -4247 -1817
rect -4199 -1831 -4195 -1817
rect -4165 -1824 -4161 -1817
rect -4235 -1860 -4231 -1841
rect -4228 -1860 -4207 -1858
rect -4231 -1863 -4207 -1860
rect -4191 -1859 -4187 -1841
rect -4157 -1852 -4153 -1834
rect -4127 -1838 -4093 -1834
rect -4121 -1844 -4117 -1838
rect -4157 -1856 -4145 -1852
rect -4191 -1863 -4164 -1859
rect -4149 -1862 -4145 -1856
rect -4103 -1861 -4099 -1854
rect -4231 -1865 -4223 -1863
rect -4251 -1870 -4247 -1865
rect -4257 -1873 -4225 -1870
rect -4207 -1882 -4203 -1876
rect -4191 -1882 -4187 -1863
rect -4149 -1866 -4119 -1862
rect -4103 -1866 -4077 -1861
rect -4207 -1886 -4187 -1882
rect -4184 -1889 -4180 -1876
rect -4103 -1869 -4099 -1866
rect -4165 -1887 -4161 -1876
rect -4121 -1880 -4117 -1874
rect -4127 -1883 -4093 -1880
rect -4210 -1894 -4176 -1889
rect -4168 -1892 -4144 -1887
rect -4012 -1910 -4007 -1278
rect -3936 -1836 -3931 -1278
rect -3496 -1386 -3462 -1382
rect -3490 -1391 -3486 -1386
rect -3472 -1391 -3468 -1386
rect -3448 -1388 -3414 -1384
rect -3442 -1394 -3438 -1388
rect -3504 -1413 -3489 -1408
rect -3481 -1415 -3477 -1401
rect -3481 -1416 -3468 -1415
rect -3459 -1416 -3440 -1412
rect -3481 -1419 -3456 -1416
rect -3472 -1420 -3456 -1419
rect -3442 -1430 -3438 -1424
rect -3490 -1434 -3486 -1430
rect -3448 -1433 -3414 -1430
rect -3496 -1437 -3462 -1434
rect -3255 -1437 -3221 -1433
rect -3370 -1447 -3336 -1443
rect -3249 -1445 -3245 -1437
rect -3364 -1455 -3360 -1447
rect -3321 -1456 -3287 -1452
rect -3315 -1462 -3311 -1456
rect -3206 -1446 -3172 -1442
rect -3200 -1452 -3196 -1446
rect -3738 -1488 -3498 -1484
rect -3830 -1504 -3796 -1500
rect -3824 -1509 -3820 -1504
rect -3806 -1509 -3802 -1504
rect -3782 -1506 -3748 -1502
rect -3776 -1512 -3772 -1506
rect -3849 -1530 -3823 -1526
rect -3849 -1577 -3843 -1530
rect -3815 -1533 -3811 -1519
rect -3758 -1530 -3754 -1522
rect -3738 -1530 -3734 -1488
rect -3726 -1495 -3692 -1491
rect -3720 -1503 -3716 -1495
rect -3677 -1504 -3643 -1500
rect -3671 -1510 -3667 -1504
rect -3815 -1534 -3802 -1533
rect -3793 -1534 -3774 -1530
rect -3758 -1534 -3719 -1530
rect -3815 -1537 -3790 -1534
rect -3758 -1537 -3754 -1534
rect -3702 -1536 -3698 -1523
rect -3653 -1527 -3649 -1520
rect -3503 -1517 -3498 -1488
rect -3346 -1488 -3342 -1475
rect -3297 -1480 -3293 -1472
rect -3286 -1476 -3248 -1472
rect -3286 -1480 -3282 -1476
rect -3231 -1478 -3227 -1465
rect -3182 -1470 -3178 -1462
rect -3155 -1470 -3150 -991
rect -2832 -1109 -2461 -1104
rect -2924 -1269 -2890 -1265
rect -2918 -1274 -2914 -1269
rect -2900 -1274 -2896 -1269
rect -2876 -1271 -2842 -1267
rect -2870 -1277 -2866 -1271
rect -2953 -1295 -2917 -1291
rect -2953 -1397 -2947 -1295
rect -2909 -1298 -2905 -1284
rect -2852 -1295 -2848 -1287
rect -2832 -1295 -2826 -1109
rect -2439 -1113 -2405 -1109
rect -2433 -1118 -2429 -1113
rect -2415 -1118 -2411 -1113
rect -2391 -1115 -2357 -1111
rect -2385 -1121 -2381 -1115
rect -2483 -1140 -2471 -1135
rect -2466 -1140 -2432 -1135
rect -2483 -1258 -2479 -1140
rect -2424 -1142 -2420 -1128
rect -2367 -1139 -2363 -1131
rect -2424 -1143 -2411 -1142
rect -2402 -1143 -2383 -1139
rect -2367 -1143 -2344 -1139
rect -2424 -1146 -2399 -1143
rect -2367 -1146 -2363 -1143
rect -2415 -1147 -2399 -1146
rect -2385 -1157 -2381 -1151
rect -2433 -1161 -2429 -1157
rect -2391 -1160 -2357 -1157
rect -2439 -1164 -2405 -1161
rect -2347 -1194 -2344 -1143
rect -2300 -1159 -2266 -1155
rect -2294 -1167 -2290 -1159
rect -2251 -1168 -2217 -1164
rect -2245 -1174 -2241 -1168
rect -2347 -1198 -2293 -1194
rect -2276 -1200 -2272 -1187
rect -2227 -1192 -2223 -1184
rect -2263 -1196 -2243 -1192
rect -2227 -1196 -2163 -1192
rect -2263 -1200 -2259 -1196
rect -2227 -1199 -2223 -1196
rect -2276 -1201 -2259 -1200
rect -2286 -1204 -2259 -1201
rect -2286 -1207 -2280 -1204
rect -2245 -1210 -2241 -1204
rect -2294 -1218 -2290 -1212
rect -2276 -1218 -2272 -1212
rect -2251 -1213 -2217 -1210
rect -2300 -1221 -2266 -1218
rect -2440 -1236 -2406 -1232
rect -2434 -1241 -2430 -1236
rect -2416 -1241 -2412 -1236
rect -2392 -1238 -2358 -1234
rect -2386 -1244 -2382 -1238
rect -2483 -1262 -2433 -1258
rect -2909 -1299 -2896 -1298
rect -2887 -1299 -2868 -1295
rect -2852 -1299 -2816 -1295
rect -2909 -1302 -2884 -1299
rect -2852 -1302 -2848 -1299
rect -2900 -1303 -2884 -1302
rect -2870 -1313 -2866 -1307
rect -2918 -1317 -2914 -1313
rect -2876 -1316 -2842 -1313
rect -2924 -1320 -2890 -1317
rect -2820 -1339 -2816 -1299
rect -2792 -1304 -2758 -1300
rect -2786 -1312 -2782 -1304
rect -2743 -1313 -2709 -1309
rect -2737 -1319 -2733 -1313
rect -2820 -1343 -2785 -1339
rect -2768 -1345 -2764 -1332
rect -2719 -1337 -2715 -1329
rect -2755 -1341 -2735 -1337
rect -2719 -1341 -2699 -1337
rect -2755 -1345 -2751 -1341
rect -2719 -1344 -2715 -1341
rect -2768 -1346 -2751 -1345
rect -2778 -1349 -2751 -1346
rect -2778 -1352 -2772 -1349
rect -2737 -1355 -2733 -1349
rect -2786 -1363 -2782 -1357
rect -2768 -1363 -2764 -1357
rect -2743 -1358 -2709 -1355
rect -2792 -1366 -2758 -1363
rect -2925 -1375 -2891 -1371
rect -2919 -1380 -2915 -1375
rect -2901 -1380 -2897 -1375
rect -2877 -1377 -2843 -1373
rect -2871 -1383 -2867 -1377
rect -2702 -1378 -2699 -1341
rect -2676 -1343 -2642 -1339
rect -2670 -1351 -2666 -1343
rect -2627 -1352 -2593 -1348
rect -2621 -1358 -2617 -1352
rect -2702 -1382 -2669 -1378
rect -2953 -1401 -2918 -1397
rect -2953 -1441 -2947 -1401
rect -2910 -1404 -2906 -1390
rect -2652 -1384 -2648 -1371
rect -2603 -1376 -2599 -1368
rect -2639 -1380 -2619 -1376
rect -2603 -1380 -2591 -1376
rect -2639 -1384 -2635 -1380
rect -2603 -1383 -2599 -1380
rect -2652 -1385 -2635 -1384
rect -2662 -1388 -2635 -1385
rect -2662 -1391 -2656 -1388
rect -2621 -1394 -2617 -1388
rect -2910 -1405 -2897 -1404
rect -2888 -1405 -2869 -1401
rect -2670 -1402 -2666 -1396
rect -2652 -1402 -2648 -1396
rect -2627 -1397 -2593 -1394
rect -2910 -1408 -2885 -1405
rect -2788 -1406 -2754 -1402
rect -2676 -1405 -2642 -1402
rect -2901 -1409 -2885 -1408
rect -2871 -1419 -2867 -1413
rect -2782 -1414 -2778 -1406
rect -2919 -1423 -2915 -1419
rect -2877 -1422 -2843 -1419
rect -2925 -1426 -2891 -1423
rect -2739 -1415 -2705 -1411
rect -2733 -1421 -2729 -1415
rect -2953 -1447 -2816 -1441
rect -3218 -1474 -3198 -1470
rect -3182 -1474 -3150 -1470
rect -2921 -1472 -2887 -1468
rect -3218 -1478 -3214 -1474
rect -3182 -1477 -3178 -1474
rect -3231 -1479 -3214 -1478
rect -3333 -1484 -3313 -1480
rect -3297 -1484 -3282 -1480
rect -3241 -1482 -3214 -1479
rect -2915 -1477 -2911 -1472
rect -2897 -1477 -2893 -1472
rect -2873 -1474 -2839 -1470
rect -3333 -1488 -3329 -1484
rect -3297 -1487 -3293 -1484
rect -3241 -1485 -3235 -1482
rect -3346 -1489 -3329 -1488
rect -3491 -1495 -3457 -1491
rect -3356 -1492 -3329 -1489
rect -3200 -1488 -3196 -1482
rect -2867 -1480 -2863 -1474
rect -3485 -1500 -3481 -1495
rect -3467 -1500 -3463 -1495
rect -3443 -1497 -3409 -1493
rect -3356 -1495 -3350 -1492
rect -3437 -1503 -3433 -1497
rect -3315 -1498 -3311 -1492
rect -3249 -1496 -3245 -1490
rect -3231 -1496 -3227 -1490
rect -3206 -1491 -3172 -1488
rect -3503 -1521 -3484 -1517
rect -3476 -1524 -3472 -1510
rect -3364 -1506 -3360 -1500
rect -3346 -1506 -3342 -1500
rect -3321 -1501 -3287 -1498
rect -3255 -1499 -3221 -1496
rect -2944 -1498 -2914 -1494
rect -3370 -1509 -3336 -1506
rect -3419 -1521 -3415 -1513
rect -3476 -1525 -3463 -1524
rect -3454 -1525 -3435 -1521
rect -3419 -1525 -3382 -1521
rect -3689 -1532 -3669 -1528
rect -3653 -1532 -3634 -1527
rect -3476 -1528 -3451 -1525
rect -3419 -1528 -3415 -1525
rect -3467 -1529 -3451 -1528
rect -3689 -1536 -3685 -1532
rect -3653 -1535 -3649 -1532
rect -3702 -1537 -3685 -1536
rect -3806 -1538 -3790 -1537
rect -3712 -1540 -3685 -1537
rect -3437 -1539 -3433 -1533
rect -3776 -1548 -3772 -1542
rect -3712 -1543 -3706 -1540
rect -3671 -1546 -3667 -1540
rect -3485 -1543 -3481 -1539
rect -3443 -1542 -3409 -1539
rect -3491 -1546 -3457 -1543
rect -3824 -1552 -3820 -1548
rect -3782 -1551 -3748 -1548
rect -3830 -1555 -3796 -1552
rect -3720 -1554 -3716 -1548
rect -3702 -1554 -3698 -1548
rect -3677 -1549 -3643 -1546
rect -3726 -1557 -3692 -1554
rect -3541 -1562 -3258 -1554
rect -3849 -1584 -3581 -1577
rect -3781 -1597 -3747 -1593
rect -3775 -1602 -3771 -1597
rect -3757 -1602 -3753 -1597
rect -3733 -1599 -3699 -1595
rect -3827 -1606 -3793 -1602
rect -3821 -1612 -3817 -1606
rect -3727 -1605 -3723 -1599
rect -3851 -1630 -3848 -1629
rect -3803 -1630 -3799 -1622
rect -3790 -1623 -3774 -1619
rect -3790 -1630 -3786 -1623
rect -3766 -1626 -3762 -1612
rect -3754 -1623 -3750 -1619
rect -3709 -1623 -3705 -1615
rect -3766 -1627 -3753 -1626
rect -3740 -1627 -3725 -1623
rect -3709 -1627 -3689 -1623
rect -3766 -1630 -3736 -1627
rect -3709 -1630 -3705 -1627
rect -3851 -1634 -3819 -1630
rect -3803 -1634 -3786 -1630
rect -3757 -1631 -3736 -1630
rect -3803 -1637 -3799 -1634
rect -3727 -1641 -3723 -1635
rect -3821 -1648 -3817 -1642
rect -3775 -1645 -3771 -1641
rect -3733 -1644 -3699 -1641
rect -3781 -1648 -3747 -1645
rect -3827 -1651 -3793 -1648
rect -3827 -1662 -3793 -1658
rect -3821 -1668 -3817 -1662
rect -3779 -1663 -3745 -1659
rect -3773 -1668 -3769 -1663
rect -3755 -1668 -3751 -1663
rect -3731 -1665 -3697 -1661
rect -3694 -1665 -3689 -1627
rect -3673 -1630 -3639 -1626
rect -3667 -1638 -3663 -1630
rect -3624 -1639 -3590 -1635
rect -3618 -1645 -3614 -1639
rect -3725 -1671 -3721 -1665
rect -3694 -1669 -3666 -1665
rect -3649 -1671 -3645 -1658
rect -3600 -1663 -3596 -1655
rect -3585 -1663 -3581 -1584
rect -3636 -1667 -3616 -1663
rect -3600 -1667 -3581 -1663
rect -3636 -1671 -3632 -1667
rect -3600 -1670 -3596 -1667
rect -3803 -1686 -3799 -1678
rect -3789 -1686 -3772 -1685
rect -3835 -1690 -3819 -1686
rect -3803 -1689 -3772 -1686
rect -3803 -1690 -3788 -1689
rect -3803 -1693 -3799 -1690
rect -3764 -1692 -3760 -1678
rect -3649 -1672 -3632 -1671
rect -3659 -1675 -3632 -1672
rect -3659 -1678 -3653 -1675
rect -3752 -1689 -3748 -1685
rect -3707 -1689 -3703 -1681
rect -3618 -1681 -3614 -1675
rect -3764 -1693 -3751 -1692
rect -3738 -1693 -3723 -1689
rect -3707 -1693 -3693 -1689
rect -3667 -1689 -3663 -1683
rect -3649 -1689 -3645 -1683
rect -3624 -1684 -3590 -1681
rect -3673 -1692 -3639 -1689
rect -3764 -1696 -3734 -1693
rect -3707 -1696 -3703 -1693
rect -3755 -1697 -3734 -1696
rect -3821 -1704 -3817 -1698
rect -3827 -1707 -3793 -1704
rect -3725 -1707 -3721 -1701
rect -3773 -1711 -3769 -1707
rect -3731 -1710 -3697 -1707
rect -3779 -1714 -3748 -1711
rect -3811 -1772 -3777 -1768
rect -3805 -1777 -3801 -1772
rect -3787 -1777 -3783 -1772
rect -3763 -1774 -3729 -1770
rect -3757 -1780 -3753 -1774
rect -3813 -1799 -3804 -1794
rect -3796 -1801 -3792 -1787
rect -3739 -1798 -3735 -1790
rect -3796 -1802 -3783 -1801
rect -3774 -1802 -3755 -1798
rect -3796 -1805 -3771 -1802
rect -3739 -1803 -3725 -1798
rect -3739 -1805 -3735 -1803
rect -3787 -1806 -3771 -1805
rect -3757 -1816 -3753 -1810
rect -3805 -1820 -3801 -1816
rect -3763 -1819 -3729 -1816
rect -3811 -1823 -3777 -1820
rect -3585 -1836 -3581 -1667
rect -3540 -1809 -3535 -1562
rect -3429 -1595 -3395 -1591
rect -3423 -1600 -3419 -1595
rect -3405 -1600 -3401 -1595
rect -3381 -1597 -3347 -1593
rect -3475 -1604 -3441 -1600
rect -3469 -1610 -3465 -1604
rect -3375 -1603 -3371 -1597
rect -3499 -1628 -3496 -1627
rect -3451 -1628 -3447 -1620
rect -3438 -1621 -3422 -1617
rect -3438 -1628 -3434 -1621
rect -3414 -1624 -3410 -1610
rect -3402 -1621 -3398 -1617
rect -3357 -1621 -3353 -1613
rect -3414 -1625 -3401 -1624
rect -3388 -1625 -3373 -1621
rect -3357 -1625 -3337 -1621
rect -3414 -1628 -3384 -1625
rect -3357 -1628 -3353 -1625
rect -3499 -1632 -3467 -1628
rect -3451 -1632 -3434 -1628
rect -3405 -1629 -3384 -1628
rect -3451 -1635 -3447 -1632
rect -3375 -1639 -3371 -1633
rect -3469 -1646 -3465 -1640
rect -3423 -1643 -3419 -1639
rect -3381 -1642 -3347 -1639
rect -3429 -1646 -3395 -1643
rect -3475 -1649 -3441 -1646
rect -3475 -1660 -3441 -1656
rect -3469 -1666 -3465 -1660
rect -3427 -1661 -3393 -1657
rect -3421 -1666 -3417 -1661
rect -3403 -1666 -3399 -1661
rect -3379 -1663 -3345 -1659
rect -3342 -1663 -3337 -1625
rect -3321 -1628 -3287 -1624
rect -3315 -1636 -3311 -1628
rect -3233 -1633 -3228 -1565
rect -3272 -1637 -3238 -1633
rect -3266 -1643 -3262 -1637
rect -3373 -1669 -3369 -1663
rect -3342 -1667 -3314 -1663
rect -3297 -1669 -3293 -1656
rect -3248 -1661 -3244 -1653
rect -3233 -1661 -3228 -1638
rect -3284 -1665 -3264 -1661
rect -3248 -1665 -3228 -1661
rect -3284 -1669 -3280 -1665
rect -3248 -1668 -3244 -1665
rect -3451 -1684 -3447 -1676
rect -3437 -1684 -3420 -1683
rect -3483 -1688 -3467 -1684
rect -3451 -1687 -3420 -1684
rect -3451 -1688 -3436 -1687
rect -3451 -1691 -3447 -1688
rect -3412 -1690 -3408 -1676
rect -3297 -1670 -3280 -1669
rect -3307 -1673 -3280 -1670
rect -3307 -1676 -3301 -1673
rect -3400 -1687 -3396 -1683
rect -3355 -1687 -3351 -1679
rect -3266 -1679 -3262 -1673
rect -3412 -1691 -3399 -1690
rect -3386 -1691 -3371 -1687
rect -3355 -1691 -3341 -1687
rect -3315 -1687 -3311 -1681
rect -3297 -1687 -3293 -1681
rect -3272 -1682 -3238 -1679
rect -3321 -1690 -3287 -1687
rect -3412 -1694 -3382 -1691
rect -3355 -1694 -3351 -1691
rect -3403 -1695 -3382 -1694
rect -3469 -1702 -3465 -1696
rect -3475 -1705 -3441 -1702
rect -3373 -1705 -3369 -1699
rect -3421 -1709 -3417 -1705
rect -3379 -1708 -3345 -1705
rect -3427 -1712 -3396 -1709
rect -3424 -1752 -3390 -1748
rect -3418 -1757 -3414 -1752
rect -3400 -1757 -3396 -1752
rect -3376 -1754 -3342 -1750
rect -3370 -1760 -3366 -1754
rect -3459 -1779 -3417 -1774
rect -3409 -1781 -3405 -1767
rect -3352 -1778 -3348 -1770
rect -3409 -1782 -3396 -1781
rect -3387 -1782 -3368 -1778
rect -3352 -1782 -3317 -1778
rect -3409 -1785 -3384 -1782
rect -3352 -1785 -3348 -1782
rect -3400 -1786 -3384 -1785
rect -3321 -1787 -3317 -1782
rect -3183 -1787 -3178 -1544
rect -2944 -1563 -2938 -1498
rect -2906 -1501 -2902 -1487
rect -2906 -1502 -2893 -1501
rect -2884 -1502 -2865 -1498
rect -2906 -1505 -2881 -1502
rect -2897 -1506 -2881 -1505
rect -2867 -1516 -2863 -1510
rect -2915 -1520 -2911 -1516
rect -2873 -1519 -2839 -1516
rect -2921 -1523 -2887 -1520
rect -2824 -1563 -2816 -1447
rect -2804 -1445 -2781 -1441
rect -2804 -1542 -2798 -1445
rect -2764 -1447 -2760 -1434
rect -2751 -1443 -2731 -1439
rect -2751 -1447 -2747 -1443
rect -2764 -1448 -2747 -1447
rect -2774 -1451 -2747 -1448
rect -2774 -1454 -2768 -1451
rect -2733 -1457 -2729 -1451
rect -2782 -1465 -2778 -1459
rect -2764 -1465 -2760 -1459
rect -2739 -1460 -2705 -1457
rect -2788 -1468 -2754 -1465
rect -2558 -1542 -2553 -1355
rect -2804 -1551 -2553 -1542
rect -2483 -1381 -2479 -1262
rect -2425 -1265 -2421 -1251
rect -2425 -1266 -2412 -1265
rect -2403 -1266 -2384 -1262
rect -2425 -1269 -2400 -1266
rect -2416 -1270 -2400 -1269
rect -2386 -1280 -2382 -1274
rect -2434 -1284 -2430 -1280
rect -2392 -1283 -2358 -1280
rect -2440 -1287 -2406 -1284
rect -2167 -1314 -2163 -1196
rect -1939 -1270 -1905 -1266
rect -2124 -1279 -2090 -1275
rect -1933 -1278 -1929 -1270
rect -1830 -1271 -1798 -1268
rect -1778 -1271 -1754 -1268
rect -1744 -1271 -1720 -1268
rect -1824 -1275 -1820 -1271
rect -2118 -1287 -2114 -1279
rect -2075 -1288 -2041 -1284
rect -2069 -1294 -2065 -1288
rect -1890 -1279 -1856 -1275
rect -1884 -1285 -1880 -1279
rect -1772 -1285 -1768 -1271
rect -1738 -1278 -1734 -1271
rect -2167 -1318 -2117 -1314
rect -2100 -1320 -2096 -1307
rect -2051 -1312 -2047 -1304
rect -2005 -1309 -1932 -1305
rect -2005 -1312 -2001 -1309
rect -1915 -1311 -1911 -1298
rect -1902 -1307 -1882 -1303
rect -1902 -1311 -1898 -1307
rect -1915 -1312 -1898 -1311
rect -2087 -1316 -2067 -1312
rect -2051 -1316 -2001 -1312
rect -1925 -1315 -1898 -1312
rect -1808 -1314 -1804 -1295
rect -1801 -1314 -1780 -1312
rect -2087 -1320 -2083 -1316
rect -2051 -1319 -2047 -1316
rect -1925 -1318 -1919 -1315
rect -2100 -1321 -2083 -1320
rect -2110 -1324 -2083 -1321
rect -1884 -1321 -1880 -1315
rect -1804 -1317 -1780 -1314
rect -1764 -1313 -1760 -1295
rect -1730 -1306 -1726 -1288
rect -1700 -1292 -1666 -1288
rect -1694 -1298 -1690 -1292
rect -1730 -1310 -1718 -1306
rect -1764 -1317 -1737 -1313
rect -1722 -1316 -1718 -1310
rect -1676 -1316 -1672 -1308
rect -1804 -1319 -1796 -1317
rect -2110 -1327 -2104 -1324
rect -2069 -1330 -2065 -1324
rect -1933 -1329 -1929 -1323
rect -1915 -1329 -1911 -1323
rect -1890 -1324 -1856 -1321
rect -1824 -1324 -1820 -1319
rect -1830 -1327 -1798 -1324
rect -2118 -1338 -2114 -1332
rect -2100 -1338 -2096 -1332
rect -2075 -1333 -2041 -1330
rect -1939 -1332 -1905 -1329
rect -1780 -1336 -1776 -1330
rect -1764 -1336 -1760 -1317
rect -1722 -1320 -1692 -1316
rect -1676 -1320 -1666 -1316
rect -2124 -1341 -2090 -1338
rect -1780 -1340 -1760 -1336
rect -1757 -1343 -1753 -1330
rect -1676 -1323 -1672 -1320
rect -1738 -1341 -1734 -1330
rect -1694 -1334 -1690 -1328
rect -1700 -1337 -1666 -1334
rect -1783 -1348 -1749 -1343
rect -1741 -1346 -1717 -1341
rect -2435 -1359 -2401 -1355
rect -2429 -1364 -2425 -1359
rect -2411 -1364 -2407 -1359
rect -2387 -1361 -2353 -1357
rect -2381 -1367 -2377 -1361
rect -2483 -1385 -2428 -1381
rect -2483 -1509 -2479 -1385
rect -2420 -1388 -2416 -1374
rect -2363 -1385 -2359 -1377
rect -2420 -1389 -2407 -1388
rect -2398 -1389 -2379 -1385
rect -2363 -1389 -2340 -1385
rect -2420 -1392 -2395 -1389
rect -2363 -1392 -2359 -1389
rect -2411 -1393 -2395 -1392
rect -2381 -1403 -2377 -1397
rect -2429 -1407 -2425 -1403
rect -2387 -1406 -2353 -1403
rect -2435 -1410 -2401 -1407
rect -2343 -1438 -2340 -1389
rect -2301 -1403 -2267 -1399
rect -2295 -1411 -2291 -1403
rect -2252 -1412 -2218 -1408
rect -2246 -1418 -2242 -1412
rect -2343 -1442 -2294 -1438
rect -2277 -1444 -2273 -1431
rect -2264 -1440 -2244 -1436
rect -2264 -1444 -2260 -1440
rect -2277 -1445 -2260 -1444
rect -2287 -1448 -2260 -1445
rect -2287 -1451 -2281 -1448
rect -2246 -1454 -2242 -1448
rect -2295 -1462 -2291 -1456
rect -2277 -1462 -2273 -1456
rect -2252 -1457 -2218 -1454
rect -2301 -1465 -2267 -1462
rect -2436 -1487 -2402 -1483
rect -2430 -1492 -2426 -1487
rect -2412 -1492 -2408 -1487
rect -2388 -1489 -2354 -1485
rect -2382 -1495 -2378 -1489
rect -2483 -1513 -2429 -1509
rect -2483 -1544 -2479 -1513
rect -2421 -1516 -2417 -1502
rect -2421 -1517 -2408 -1516
rect -2399 -1517 -2380 -1513
rect -2421 -1520 -2396 -1517
rect -2412 -1521 -2396 -1520
rect -2382 -1531 -2378 -1525
rect -2430 -1535 -2426 -1531
rect -2388 -1534 -2354 -1531
rect -2436 -1538 -2402 -1535
rect -2483 -1550 -1993 -1544
rect -2944 -1568 -2668 -1563
rect -2868 -1595 -2834 -1591
rect -2862 -1600 -2858 -1595
rect -2844 -1600 -2840 -1595
rect -2820 -1597 -2786 -1593
rect -2914 -1604 -2880 -1600
rect -2908 -1610 -2904 -1604
rect -2814 -1603 -2810 -1597
rect -2938 -1632 -2906 -1627
rect -2890 -1628 -2886 -1620
rect -2877 -1621 -2861 -1617
rect -2877 -1628 -2873 -1621
rect -2853 -1624 -2849 -1610
rect -2841 -1621 -2837 -1617
rect -2796 -1621 -2792 -1613
rect -2853 -1625 -2840 -1624
rect -2827 -1625 -2812 -1621
rect -2796 -1625 -2776 -1621
rect -2853 -1628 -2823 -1625
rect -2796 -1628 -2792 -1625
rect -2890 -1632 -2873 -1628
rect -2844 -1629 -2823 -1628
rect -3370 -1796 -3366 -1790
rect -3321 -1791 -3178 -1787
rect -2890 -1635 -2886 -1632
rect -3418 -1800 -3414 -1796
rect -3376 -1799 -3342 -1796
rect -3424 -1803 -3390 -1800
rect -3321 -1809 -3317 -1791
rect -3540 -1814 -3317 -1809
rect -3936 -1840 -3581 -1836
rect -3139 -1910 -3134 -1638
rect -2814 -1639 -2810 -1633
rect -2908 -1646 -2904 -1640
rect -2862 -1643 -2858 -1639
rect -2820 -1642 -2786 -1639
rect -2868 -1646 -2834 -1643
rect -2914 -1649 -2880 -1646
rect -2914 -1660 -2880 -1656
rect -2908 -1666 -2904 -1660
rect -2866 -1661 -2832 -1657
rect -2860 -1666 -2856 -1661
rect -2842 -1666 -2838 -1661
rect -2818 -1663 -2784 -1659
rect -2781 -1663 -2776 -1625
rect -2760 -1628 -2726 -1624
rect -2754 -1636 -2750 -1628
rect -2711 -1637 -2677 -1633
rect -2705 -1643 -2701 -1637
rect -2812 -1669 -2808 -1663
rect -2781 -1667 -2753 -1663
rect -2736 -1669 -2732 -1656
rect -2687 -1661 -2683 -1653
rect -2673 -1660 -2668 -1568
rect -2723 -1665 -2703 -1661
rect -2687 -1665 -2673 -1661
rect -2723 -1669 -2719 -1665
rect -2687 -1668 -2683 -1665
rect -2890 -1684 -2886 -1676
rect -2876 -1684 -2859 -1683
rect -2922 -1688 -2906 -1684
rect -2890 -1687 -2859 -1684
rect -2890 -1688 -2875 -1687
rect -2890 -1691 -2886 -1688
rect -2851 -1690 -2847 -1676
rect -2736 -1670 -2719 -1669
rect -2746 -1673 -2719 -1670
rect -2746 -1676 -2740 -1673
rect -2839 -1687 -2835 -1683
rect -2794 -1687 -2790 -1679
rect -2705 -1679 -2701 -1673
rect -2851 -1691 -2838 -1690
rect -2825 -1691 -2810 -1687
rect -2794 -1691 -2780 -1687
rect -2754 -1687 -2750 -1681
rect -2736 -1687 -2732 -1681
rect -2711 -1682 -2677 -1679
rect -2760 -1690 -2726 -1687
rect -2851 -1694 -2821 -1691
rect -2794 -1694 -2790 -1691
rect -2842 -1695 -2821 -1694
rect -2908 -1702 -2904 -1696
rect -2914 -1705 -2880 -1702
rect -2812 -1705 -2808 -1699
rect -2860 -1709 -2856 -1705
rect -2818 -1708 -2784 -1705
rect -2866 -1712 -2835 -1709
rect -2874 -1751 -2840 -1747
rect -2868 -1756 -2864 -1751
rect -2850 -1756 -2846 -1751
rect -2826 -1753 -2792 -1749
rect -2820 -1759 -2816 -1753
rect -2898 -1778 -2867 -1773
rect -2859 -1780 -2855 -1766
rect -2802 -1777 -2798 -1769
rect -2608 -1777 -2600 -1551
rect -2193 -1576 -2159 -1572
rect -2187 -1581 -2183 -1576
rect -2169 -1581 -2165 -1576
rect -2145 -1578 -2111 -1574
rect -2239 -1585 -2205 -1581
rect -2233 -1591 -2229 -1585
rect -2139 -1584 -2135 -1578
rect -2263 -1609 -2260 -1608
rect -2215 -1609 -2211 -1601
rect -2202 -1602 -2186 -1598
rect -2202 -1609 -2198 -1602
rect -2178 -1605 -2174 -1591
rect -2166 -1602 -2162 -1598
rect -2121 -1602 -2117 -1594
rect -2178 -1606 -2165 -1605
rect -2152 -1606 -2137 -1602
rect -2121 -1606 -2101 -1602
rect -2178 -1609 -2148 -1606
rect -2121 -1609 -2117 -1606
rect -2263 -1613 -2231 -1609
rect -2215 -1613 -2198 -1609
rect -2169 -1610 -2148 -1609
rect -2215 -1616 -2211 -1613
rect -2139 -1620 -2135 -1614
rect -2233 -1627 -2229 -1621
rect -2187 -1624 -2183 -1620
rect -2145 -1623 -2111 -1620
rect -2193 -1627 -2159 -1624
rect -2239 -1630 -2205 -1627
rect -2239 -1641 -2205 -1637
rect -2233 -1647 -2229 -1641
rect -2191 -1642 -2157 -1638
rect -2185 -1647 -2181 -1642
rect -2167 -1647 -2163 -1642
rect -2143 -1644 -2109 -1640
rect -2106 -1644 -2101 -1606
rect -2085 -1609 -2051 -1605
rect -2079 -1617 -2075 -1609
rect -2036 -1618 -2002 -1614
rect -2030 -1624 -2026 -1618
rect -2137 -1650 -2133 -1644
rect -2106 -1648 -2078 -1644
rect -2061 -1650 -2057 -1637
rect -2012 -1642 -2008 -1634
rect -1997 -1642 -1993 -1550
rect -2048 -1646 -2028 -1642
rect -2012 -1646 -1993 -1642
rect -2048 -1650 -2044 -1646
rect -2012 -1649 -2008 -1646
rect -2215 -1665 -2211 -1657
rect -2201 -1665 -2184 -1664
rect -2247 -1669 -2231 -1665
rect -2215 -1668 -2184 -1665
rect -2215 -1669 -2200 -1668
rect -2254 -1743 -2247 -1669
rect -2215 -1672 -2211 -1669
rect -2176 -1671 -2172 -1657
rect -2061 -1651 -2044 -1650
rect -2071 -1654 -2044 -1651
rect -2071 -1657 -2065 -1654
rect -2030 -1660 -2026 -1654
rect -2164 -1668 -2160 -1664
rect -2079 -1668 -2075 -1662
rect -2061 -1668 -2057 -1662
rect -2036 -1663 -2002 -1660
rect -2176 -1672 -2163 -1671
rect -2150 -1672 -2135 -1668
rect -2085 -1671 -2051 -1668
rect -2176 -1675 -2146 -1672
rect -2167 -1676 -2146 -1675
rect -2233 -1683 -2229 -1677
rect -2239 -1686 -2205 -1683
rect -2137 -1686 -2133 -1680
rect -2185 -1690 -2181 -1686
rect -2143 -1689 -2109 -1686
rect -2191 -1693 -2160 -1690
rect -2204 -1721 -2170 -1717
rect -2198 -1726 -2194 -1721
rect -2180 -1726 -2176 -1721
rect -2156 -1723 -2122 -1719
rect -2150 -1729 -2146 -1723
rect -2254 -1747 -2197 -1743
rect -2189 -1750 -2185 -1736
rect -2189 -1751 -2176 -1750
rect -2167 -1751 -2148 -1747
rect -2189 -1754 -2164 -1751
rect -2180 -1755 -2164 -1754
rect -2150 -1765 -2146 -1759
rect -2198 -1769 -2194 -1765
rect -2156 -1768 -2122 -1765
rect -2204 -1772 -2170 -1769
rect -2859 -1781 -2846 -1780
rect -2837 -1781 -2818 -1777
rect -2802 -1781 -2600 -1777
rect -2859 -1784 -2834 -1781
rect -2802 -1784 -2798 -1781
rect -2850 -1785 -2834 -1784
rect -2820 -1795 -2816 -1789
rect -2868 -1799 -2864 -1795
rect -2826 -1798 -2792 -1795
rect -1954 -1798 -1922 -1795
rect -1902 -1798 -1878 -1795
rect -1868 -1798 -1844 -1795
rect -2874 -1802 -2840 -1799
rect -1948 -1802 -1944 -1798
rect -2271 -1805 -2239 -1802
rect -2219 -1805 -2195 -1802
rect -2185 -1805 -2161 -1802
rect -2265 -1809 -2261 -1805
rect -2720 -1816 -2688 -1813
rect -2668 -1816 -2644 -1813
rect -2634 -1816 -2610 -1813
rect -2958 -1820 -2926 -1817
rect -2906 -1820 -2882 -1817
rect -2872 -1820 -2848 -1817
rect -2714 -1820 -2710 -1816
rect -2952 -1824 -2948 -1820
rect -2900 -1834 -2896 -1820
rect -2866 -1827 -2862 -1820
rect -2936 -1863 -2932 -1844
rect -2929 -1863 -2908 -1861
rect -2932 -1866 -2908 -1863
rect -2892 -1862 -2888 -1844
rect -2858 -1855 -2854 -1837
rect -2828 -1841 -2794 -1837
rect -2662 -1830 -2658 -1816
rect -2628 -1823 -2624 -1816
rect -2213 -1819 -2209 -1805
rect -2179 -1812 -2175 -1805
rect -1896 -1812 -1892 -1798
rect -1862 -1805 -1858 -1798
rect -2822 -1847 -2818 -1841
rect -2858 -1859 -2846 -1855
rect -2892 -1866 -2865 -1862
rect -2850 -1865 -2846 -1859
rect -2804 -1864 -2800 -1857
rect -2698 -1859 -2694 -1840
rect -2691 -1859 -2670 -1857
rect -2694 -1862 -2670 -1859
rect -2654 -1858 -2650 -1840
rect -2620 -1851 -2616 -1833
rect -2590 -1837 -2556 -1833
rect -2584 -1843 -2580 -1837
rect -2620 -1855 -2608 -1851
rect -2249 -1848 -2245 -1829
rect -2242 -1848 -2221 -1846
rect -2654 -1862 -2627 -1858
rect -2612 -1861 -2608 -1855
rect -2566 -1860 -2562 -1853
rect -2245 -1851 -2221 -1848
rect -2205 -1847 -2201 -1829
rect -2171 -1840 -2167 -1822
rect -2141 -1826 -2107 -1822
rect -2135 -1832 -2131 -1826
rect -2171 -1844 -2159 -1840
rect -1932 -1841 -1928 -1822
rect -1925 -1841 -1904 -1839
rect -2205 -1851 -2178 -1847
rect -2163 -1850 -2159 -1844
rect -2117 -1849 -2113 -1842
rect -1928 -1844 -1904 -1841
rect -1888 -1840 -1884 -1822
rect -1854 -1833 -1850 -1815
rect -1824 -1819 -1790 -1815
rect -1818 -1825 -1814 -1819
rect -1854 -1837 -1842 -1833
rect -1888 -1844 -1861 -1840
rect -1846 -1843 -1842 -1837
rect -1800 -1842 -1796 -1835
rect -1928 -1846 -1920 -1844
rect -2245 -1853 -2237 -1851
rect -2265 -1858 -2261 -1853
rect -2694 -1864 -2686 -1862
rect -2932 -1868 -2924 -1866
rect -2952 -1873 -2948 -1868
rect -2958 -1876 -2926 -1873
rect -2908 -1885 -2904 -1879
rect -2892 -1885 -2888 -1866
rect -2850 -1869 -2820 -1865
rect -2804 -1869 -2791 -1864
rect -2714 -1869 -2710 -1864
rect -2908 -1889 -2888 -1885
rect -2885 -1892 -2881 -1879
rect -2804 -1872 -2800 -1869
rect -2720 -1872 -2688 -1869
rect -2866 -1890 -2862 -1879
rect -2822 -1883 -2818 -1877
rect -2670 -1881 -2666 -1875
rect -2654 -1881 -2650 -1862
rect -2612 -1865 -2582 -1861
rect -2566 -1865 -2552 -1860
rect -2271 -1861 -2239 -1858
rect -2828 -1886 -2794 -1883
rect -2670 -1885 -2650 -1881
rect -2647 -1888 -2643 -1875
rect -2566 -1868 -2562 -1865
rect -2221 -1870 -2217 -1864
rect -2205 -1870 -2201 -1851
rect -2163 -1854 -2133 -1850
rect -2117 -1854 -2105 -1849
rect -1948 -1851 -1944 -1846
rect -1954 -1854 -1922 -1851
rect -2628 -1886 -2624 -1875
rect -2584 -1879 -2580 -1873
rect -2221 -1874 -2201 -1870
rect -2198 -1877 -2194 -1864
rect -2117 -1857 -2113 -1854
rect -2179 -1875 -2175 -1864
rect -2135 -1868 -2131 -1862
rect -1904 -1863 -1900 -1857
rect -1888 -1863 -1884 -1844
rect -1846 -1847 -1816 -1843
rect -1800 -1847 -1781 -1842
rect -1904 -1867 -1884 -1863
rect -2141 -1871 -2107 -1868
rect -1881 -1870 -1877 -1857
rect -1800 -1850 -1796 -1847
rect -1862 -1868 -1858 -1857
rect -1818 -1861 -1814 -1855
rect -1824 -1864 -1790 -1861
rect -1907 -1875 -1873 -1870
rect -1865 -1873 -1841 -1868
rect -2590 -1882 -2556 -1879
rect -2224 -1882 -2190 -1877
rect -2182 -1880 -2158 -1875
rect -2911 -1897 -2877 -1892
rect -2869 -1895 -2845 -1890
rect -2673 -1893 -2639 -1888
rect -2631 -1891 -2607 -1886
rect -4012 -1917 -3134 -1910
rect -3334 -1969 -3302 -1966
rect -3282 -1969 -3258 -1966
rect -3248 -1969 -3224 -1966
rect -3328 -1973 -3324 -1969
rect -3633 -1978 -3601 -1975
rect -3581 -1978 -3557 -1975
rect -3547 -1978 -3523 -1975
rect -3627 -1982 -3623 -1978
rect -3575 -1992 -3571 -1978
rect -3541 -1985 -3537 -1978
rect -3276 -1983 -3272 -1969
rect -3242 -1976 -3238 -1969
rect -3611 -2021 -3607 -2002
rect -3604 -2021 -3583 -2019
rect -3607 -2024 -3583 -2021
rect -3567 -2020 -3563 -2002
rect -3533 -2013 -3529 -1995
rect -3503 -1999 -3469 -1995
rect -3497 -2005 -3493 -1999
rect -3533 -2017 -3521 -2013
rect -3312 -2012 -3308 -1993
rect -3305 -2012 -3284 -2010
rect -3567 -2024 -3540 -2020
rect -3525 -2023 -3521 -2017
rect -3479 -2022 -3475 -2015
rect -3308 -2015 -3284 -2012
rect -3268 -2011 -3264 -1993
rect -3234 -2004 -3230 -1986
rect -3204 -1990 -3170 -1986
rect -3198 -1996 -3194 -1990
rect -3234 -2008 -3222 -2004
rect -3268 -2015 -3241 -2011
rect -3226 -2014 -3222 -2008
rect -3180 -2013 -3176 -2006
rect -3166 -2013 -3161 -1932
rect -3308 -2017 -3300 -2015
rect -3328 -2022 -3324 -2017
rect -3607 -2026 -3599 -2024
rect -3627 -2031 -3623 -2026
rect -3633 -2034 -3601 -2031
rect -3583 -2043 -3579 -2037
rect -3567 -2043 -3563 -2024
rect -3525 -2027 -3495 -2023
rect -3479 -2027 -3456 -2022
rect -3334 -2025 -3302 -2022
rect -3583 -2047 -3563 -2043
rect -3560 -2050 -3556 -2037
rect -3479 -2030 -3475 -2027
rect -3284 -2034 -3280 -2028
rect -3268 -2034 -3264 -2015
rect -3226 -2018 -3196 -2014
rect -3180 -2018 -3161 -2013
rect -3541 -2048 -3537 -2037
rect -3497 -2041 -3493 -2035
rect -3284 -2038 -3264 -2034
rect -3261 -2041 -3257 -2028
rect -3180 -2021 -3176 -2018
rect -3242 -2039 -3238 -2028
rect -3198 -2032 -3194 -2026
rect -3204 -2035 -3170 -2032
rect -3503 -2044 -3469 -2041
rect -3287 -2046 -3253 -2041
rect -3245 -2044 -3221 -2039
rect -3586 -2055 -3552 -2050
rect -3544 -2053 -3520 -2048
<< m2contact >>
rect -2574 -759 -2567 -752
rect -3295 -783 -3288 -778
rect -3309 -798 -3304 -793
rect -3203 -788 -3198 -783
rect -3036 -831 -3029 -826
rect -3295 -854 -3288 -849
rect -3201 -854 -3196 -849
rect -3146 -857 -3141 -852
rect -2588 -772 -2583 -767
rect -2482 -762 -2477 -757
rect -1966 -754 -1961 -749
rect -1860 -744 -1855 -739
rect -1687 -787 -1681 -782
rect -2311 -805 -2306 -800
rect -2574 -828 -2567 -823
rect -1952 -810 -1945 -805
rect -2480 -828 -2475 -823
rect -1858 -810 -1853 -805
rect -2425 -831 -2420 -826
rect -3936 -1032 -3931 -1027
rect -3854 -1044 -3849 -1039
rect -3748 -1034 -3743 -1029
rect -3552 -1077 -3543 -1072
rect -3840 -1100 -3833 -1095
rect -3746 -1100 -3741 -1095
rect -3691 -1103 -3686 -1098
rect -4131 -1364 -4126 -1359
rect -4095 -1675 -4090 -1670
rect -4082 -1861 -4077 -1856
rect -3509 -1413 -3504 -1408
rect -2461 -1109 -2456 -1104
rect -2471 -1140 -2466 -1135
rect -2558 -1355 -2553 -1350
rect -2591 -1380 -2586 -1375
rect -3388 -1521 -3382 -1516
rect -3634 -1532 -3629 -1527
rect -3183 -1544 -3178 -1539
rect -3266 -1554 -3258 -1547
rect -3856 -1634 -3851 -1629
rect -3750 -1624 -3745 -1619
rect -3842 -1690 -3835 -1685
rect -3748 -1690 -3743 -1685
rect -3693 -1693 -3688 -1688
rect -3818 -1799 -3813 -1794
rect -3725 -1803 -3720 -1798
rect -3240 -1572 -3233 -1565
rect -3504 -1632 -3499 -1627
rect -3398 -1622 -3393 -1617
rect -3233 -1638 -3228 -1633
rect -3490 -1688 -3483 -1683
rect -3396 -1688 -3391 -1683
rect -3341 -1691 -3336 -1686
rect -3464 -1779 -3459 -1774
rect -2945 -1632 -2938 -1627
rect -2837 -1622 -2832 -1617
rect -3139 -1638 -3134 -1633
rect -2673 -1665 -2668 -1660
rect -2929 -1688 -2922 -1683
rect -2835 -1688 -2830 -1683
rect -2780 -1691 -2775 -1686
rect -2903 -1778 -2898 -1773
rect -2268 -1613 -2263 -1608
rect -2162 -1603 -2157 -1598
rect -2254 -1669 -2247 -1664
rect -2160 -1669 -2155 -1664
rect -2791 -1869 -2786 -1864
rect -2552 -1865 -2547 -1860
rect -2105 -1854 -2100 -1849
rect -1781 -1847 -1775 -1842
rect -3166 -1932 -3161 -1927
rect -3456 -2027 -3451 -2022
<< metal2 >>
rect -1687 -532 -1661 -528
rect -2311 -553 -2291 -549
rect -3310 -562 -3290 -558
rect -3868 -603 -3850 -599
rect -3868 -658 -3863 -603
rect -3868 -667 -3543 -658
rect -3840 -999 -3739 -995
rect -3840 -1027 -3833 -999
rect -3931 -1032 -3833 -1027
rect -3854 -1125 -3849 -1044
rect -3840 -1095 -3833 -1032
rect -3743 -1034 -3739 -999
rect -3552 -1072 -3543 -667
rect -3310 -672 -3305 -562
rect -3310 -678 -3029 -672
rect -3295 -753 -3194 -749
rect -3295 -778 -3288 -753
rect -3309 -865 -3304 -798
rect -3295 -849 -3288 -783
rect -3198 -788 -3194 -753
rect -3036 -826 -3029 -678
rect -2574 -727 -2473 -723
rect -2574 -752 -2567 -727
rect -3111 -833 -3105 -829
rect -3146 -836 -3108 -833
rect -3309 -879 -3304 -875
rect -3201 -879 -3196 -854
rect -3146 -852 -3141 -836
rect -2588 -853 -2583 -772
rect -2574 -823 -2567 -759
rect -2477 -762 -2473 -727
rect -2311 -800 -2306 -553
rect -1952 -709 -1851 -705
rect -1952 -716 -1945 -709
rect -1969 -754 -1966 -749
rect -1969 -766 -1961 -754
rect -2391 -807 -2388 -803
rect -2026 -771 -1961 -766
rect -2425 -810 -2388 -807
rect -2480 -853 -2475 -828
rect -2425 -826 -2420 -810
rect -2588 -859 -2536 -853
rect -2530 -859 -2475 -853
rect -2026 -867 -2022 -771
rect -1969 -835 -1961 -771
rect -1952 -805 -1945 -721
rect -1855 -744 -1851 -709
rect -1687 -782 -1681 -532
rect -1769 -789 -1766 -785
rect -1803 -792 -1766 -789
rect -1858 -835 -1853 -810
rect -1817 -809 -1813 -801
rect -1803 -809 -1798 -792
rect -1817 -813 -1798 -809
rect -1817 -816 -1813 -813
rect -1969 -840 -1853 -835
rect -3309 -885 -3196 -879
rect -2347 -871 -2022 -867
rect -3656 -1079 -3650 -1075
rect -3691 -1082 -3653 -1079
rect -3746 -1125 -3741 -1100
rect -3691 -1098 -3686 -1082
rect -2347 -1087 -2344 -871
rect -2471 -1091 -2344 -1087
rect -3848 -1131 -3741 -1125
rect -2471 -1135 -2466 -1091
rect -2456 -1109 -2398 -1104
rect -2402 -1135 -2398 -1109
rect -2412 -1139 -2398 -1135
rect -2286 -1198 -2283 -1194
rect -2347 -1201 -2283 -1198
rect -2811 -1232 -2399 -1228
rect -2811 -1343 -2808 -1232
rect -2403 -1258 -2399 -1232
rect -2413 -1262 -2399 -1258
rect -2368 -1263 -2364 -1254
rect -2347 -1263 -2344 -1201
rect -2368 -1266 -2344 -1263
rect -2368 -1269 -2364 -1266
rect -1866 -1303 -1862 -1295
rect -1925 -1309 -1922 -1305
rect -1978 -1312 -1922 -1309
rect -1866 -1307 -1823 -1303
rect -1866 -1310 -1862 -1307
rect -2110 -1318 -2107 -1314
rect -2139 -1321 -2107 -1318
rect -2778 -1343 -2775 -1339
rect -2834 -1346 -2775 -1343
rect -4316 -1351 -4303 -1347
rect -4131 -1359 -4126 -1354
rect -3458 -1382 -3395 -1378
rect -3458 -1408 -3454 -1382
rect -3759 -1413 -3509 -1408
rect -3469 -1412 -3454 -1408
rect -3759 -1484 -3754 -1413
rect -3400 -1483 -3395 -1382
rect -2853 -1402 -2849 -1393
rect -2834 -1402 -2830 -1346
rect -2553 -1355 -2394 -1350
rect -2591 -1375 -2586 -1369
rect -2662 -1382 -2659 -1378
rect -2398 -1381 -2394 -1355
rect -2853 -1406 -2830 -1402
rect -2700 -1385 -2659 -1382
rect -2408 -1385 -2394 -1381
rect -2853 -1408 -2849 -1406
rect -2715 -1439 -2711 -1431
rect -2700 -1439 -2696 -1385
rect -2228 -1436 -2224 -1428
rect -2139 -1436 -2134 -1321
rect -2774 -1445 -2771 -1441
rect -2798 -1448 -2771 -1445
rect -2715 -1443 -2696 -1439
rect -2287 -1442 -2284 -1438
rect -2715 -1446 -2711 -1443
rect -2343 -1445 -2284 -1442
rect -2228 -1440 -2134 -1436
rect -2228 -1443 -2224 -1440
rect -2987 -1467 -2879 -1463
rect -3241 -1476 -3238 -1472
rect -3266 -1479 -3238 -1476
rect -3920 -1489 -3738 -1484
rect -4287 -1662 -4269 -1658
rect -4090 -1675 -4085 -1670
rect -3920 -1831 -3914 -1489
rect -3742 -1534 -3738 -1489
rect -3454 -1487 -3395 -1483
rect -3356 -1486 -3353 -1482
rect -3454 -1517 -3450 -1487
rect -3464 -1521 -3450 -1517
rect -3634 -1527 -3629 -1522
rect -3712 -1534 -3709 -1530
rect -3742 -1537 -3709 -1534
rect -3400 -1565 -3395 -1487
rect -3388 -1489 -3353 -1486
rect -3388 -1509 -3382 -1489
rect -3388 -1516 -3382 -1514
rect -3266 -1547 -3258 -1479
rect -2987 -1514 -2981 -1467
rect -2883 -1494 -2879 -1467
rect -2798 -1479 -2793 -1448
rect -2798 -1483 -2395 -1479
rect -2894 -1498 -2879 -1494
rect -2849 -1498 -2845 -1490
rect -2798 -1498 -2793 -1483
rect -2849 -1502 -2793 -1498
rect -2849 -1505 -2845 -1502
rect -2399 -1509 -2395 -1483
rect -2409 -1513 -2395 -1509
rect -3183 -1519 -2981 -1514
rect -2364 -1514 -2360 -1505
rect -2343 -1514 -2340 -1445
rect -2364 -1517 -2340 -1514
rect -3183 -1539 -3178 -1519
rect -2364 -1520 -2360 -1517
rect -3400 -1572 -3240 -1565
rect -2254 -1568 -2153 -1565
rect -2254 -1582 -2247 -1568
rect -3842 -1589 -3741 -1586
rect -3842 -1607 -3835 -1589
rect -3879 -1615 -3835 -1607
rect -3879 -1760 -3871 -1615
rect -3858 -1634 -3856 -1629
rect -3858 -1670 -3851 -1634
rect -3858 -1715 -3851 -1675
rect -3842 -1685 -3835 -1615
rect -3745 -1624 -3741 -1589
rect -3490 -1587 -3389 -1584
rect -3490 -1616 -3483 -1587
rect -3530 -1622 -3483 -1616
rect -3393 -1622 -3389 -1587
rect -2929 -1587 -2828 -1584
rect -2929 -1616 -2922 -1587
rect -2972 -1620 -2922 -1616
rect -3658 -1669 -3652 -1665
rect -3693 -1672 -3655 -1669
rect -3748 -1715 -3743 -1690
rect -3693 -1688 -3688 -1672
rect -3858 -1721 -3743 -1715
rect -3879 -1794 -3871 -1766
rect -3775 -1794 -3770 -1721
rect -3530 -1774 -3524 -1622
rect -3506 -1632 -3504 -1627
rect -3506 -1713 -3499 -1632
rect -3490 -1683 -3483 -1622
rect -3228 -1638 -3139 -1633
rect -3307 -1667 -3304 -1663
rect -3341 -1670 -3304 -1667
rect -3396 -1713 -3391 -1688
rect -3341 -1686 -3336 -1670
rect -2972 -1680 -2967 -1620
rect -3506 -1719 -3391 -1713
rect -3429 -1727 -3424 -1719
rect -3429 -1740 -3424 -1732
rect -3429 -1744 -3382 -1740
rect -3386 -1774 -3382 -1744
rect -3530 -1779 -3516 -1774
rect -3509 -1779 -3464 -1774
rect -3397 -1778 -3382 -1774
rect -2972 -1773 -2967 -1686
rect -2945 -1713 -2938 -1632
rect -2929 -1683 -2922 -1620
rect -2832 -1622 -2828 -1587
rect -2270 -1613 -2268 -1608
rect -2746 -1667 -2743 -1663
rect -2668 -1665 -2663 -1660
rect -2780 -1670 -2743 -1667
rect -2835 -1713 -2830 -1688
rect -2780 -1686 -2775 -1670
rect -2270 -1694 -2263 -1613
rect -2254 -1664 -2247 -1591
rect -2157 -1603 -2153 -1568
rect -2071 -1648 -2068 -1644
rect -2105 -1651 -2068 -1648
rect -2160 -1694 -2155 -1669
rect -2119 -1668 -2115 -1660
rect -2105 -1668 -2100 -1651
rect -2119 -1672 -2100 -1668
rect -2119 -1675 -2115 -1672
rect -2270 -1700 -2155 -1694
rect -2945 -1719 -2830 -1713
rect -2167 -1711 -2162 -1700
rect -2837 -1734 -2832 -1719
rect -2837 -1773 -2832 -1739
rect -2167 -1743 -2162 -1716
rect -2177 -1747 -2162 -1743
rect -2132 -1747 -2128 -1739
rect -1978 -1747 -1974 -1312
rect -2132 -1751 -1974 -1747
rect -2132 -1754 -2128 -1751
rect -2972 -1778 -2903 -1773
rect -2847 -1777 -2832 -1773
rect -3879 -1799 -3818 -1794
rect -3784 -1798 -3770 -1794
rect -3725 -1831 -3720 -1803
rect -3920 -1836 -3720 -1831
rect -1965 -1834 -1947 -1830
rect -2282 -1841 -2264 -1837
rect -1781 -1842 -1775 -1837
rect -4268 -1853 -4250 -1849
rect -4082 -1856 -4077 -1851
rect -2731 -1852 -2713 -1848
rect -2969 -1856 -2951 -1852
rect -2552 -1860 -2547 -1855
rect -2105 -1859 -2100 -1854
rect -2791 -1874 -2786 -1869
rect -3171 -1932 -3166 -1927
rect -3345 -2005 -3327 -2001
rect -3644 -2014 -3626 -2010
rect -3456 -2022 -3451 -2017
<< m3contact >>
rect -3309 -875 -3304 -865
rect -1952 -721 -1945 -716
rect -2536 -859 -2530 -853
rect -3854 -1131 -3848 -1125
rect -4131 -1354 -4126 -1349
rect -2591 -1369 -2586 -1363
rect -4085 -1675 -4080 -1670
rect -3634 -1522 -3629 -1517
rect -3388 -1514 -3382 -1509
rect -3858 -1675 -3851 -1670
rect -3879 -1766 -3871 -1760
rect -2972 -1686 -2967 -1680
rect -3429 -1732 -3424 -1727
rect -3516 -1779 -3509 -1774
rect -2254 -1591 -2247 -1582
rect -2663 -1665 -2658 -1660
rect -2167 -1716 -2162 -1711
rect -2837 -1739 -2832 -1734
rect -1781 -1837 -1775 -1832
rect -4082 -1851 -4077 -1846
rect -2552 -1855 -2547 -1850
rect -2105 -1864 -2100 -1859
rect -2791 -1879 -2786 -1874
rect -3176 -1932 -3171 -1927
rect -3456 -2017 -3451 -2012
<< metal3 >>
rect -2257 -448 -1282 -445
rect -2257 -503 -2253 -448
rect -3816 -508 -2253 -503
rect -3816 -547 -3811 -508
rect -4250 -553 -3811 -547
rect -3256 -509 -2253 -508
rect -3256 -519 -3252 -509
rect -2257 -510 -2253 -509
rect -1627 -489 -1623 -448
rect -1627 -493 -1549 -489
rect -2257 -514 -2179 -510
rect -3256 -523 -3178 -519
rect -4250 -1308 -4243 -553
rect -3816 -560 -3812 -553
rect -3256 -559 -3252 -523
rect -3816 -564 -3738 -560
rect -3263 -563 -3238 -559
rect -3182 -563 -3178 -523
rect -2257 -550 -2253 -514
rect -2264 -554 -2239 -550
rect -2183 -554 -2179 -514
rect -1627 -529 -1623 -493
rect -1634 -533 -1609 -529
rect -1553 -533 -1549 -493
rect -3816 -600 -3812 -564
rect -3823 -604 -3798 -600
rect -3742 -604 -3738 -564
rect -2607 -721 -1952 -716
rect -3379 -875 -3309 -865
rect -3891 -1131 -3854 -1125
rect -3379 -1126 -3368 -875
rect -2607 -878 -2602 -721
rect -2607 -885 -2586 -878
rect -3891 -1271 -3886 -1131
rect -4131 -1278 -3886 -1271
rect -4269 -1312 -4191 -1308
rect -4269 -1348 -4265 -1312
rect -4276 -1352 -4251 -1348
rect -4195 -1352 -4191 -1312
rect -4131 -1349 -4126 -1278
rect -4269 -1409 -4265 -1352
rect -4269 -1413 -4231 -1409
rect -4235 -1588 -4231 -1413
rect -3891 -1469 -3886 -1278
rect -3634 -1133 -3368 -1126
rect -3891 -1475 -3789 -1469
rect -3794 -1526 -3789 -1475
rect -3634 -1517 -3629 -1133
rect -2980 -1263 -2882 -1258
rect -2980 -1372 -2975 -1263
rect -2886 -1291 -2882 -1263
rect -2897 -1295 -2882 -1291
rect -2591 -1363 -2586 -885
rect -3395 -1376 -2975 -1372
rect -2961 -1370 -2885 -1365
rect -3424 -1412 -3420 -1404
rect -3395 -1412 -3391 -1376
rect -3424 -1416 -3391 -1412
rect -3424 -1419 -3420 -1416
rect -3395 -1482 -3391 -1416
rect -3395 -1486 -3363 -1482
rect -2961 -1509 -2956 -1370
rect -2890 -1397 -2885 -1370
rect -2898 -1401 -2885 -1397
rect -3382 -1514 -2956 -1509
rect -3803 -1530 -3789 -1526
rect -4404 -1592 -4231 -1588
rect -4404 -1767 -4398 -1592
rect -4235 -1619 -4231 -1592
rect -4235 -1623 -4157 -1619
rect -4235 -1659 -4231 -1623
rect -4242 -1663 -4217 -1659
rect -4161 -1663 -4157 -1623
rect -2536 -1660 -2530 -859
rect -1287 -1264 -1282 -448
rect -1789 -1268 -1282 -1264
rect -1789 -1304 -1785 -1268
rect -1796 -1308 -1771 -1304
rect -1715 -1308 -1711 -1268
rect -2658 -1665 -2530 -1660
rect -2324 -1591 -2254 -1582
rect -4080 -1675 -3858 -1670
rect -2978 -1686 -2972 -1680
rect -3424 -1732 -3292 -1727
rect -4082 -1766 -3879 -1760
rect -4404 -1772 -4212 -1767
rect -4321 -2086 -4315 -1772
rect -4216 -1810 -4212 -1772
rect -4216 -1814 -4138 -1810
rect -4216 -1850 -4212 -1814
rect -4223 -1854 -4198 -1850
rect -4142 -1854 -4138 -1814
rect -4082 -1846 -4077 -1766
rect -3516 -1949 -3509 -1779
rect -3297 -1927 -3292 -1732
rect -2978 -1909 -2973 -1686
rect -2832 -1739 -2547 -1734
rect -2758 -1809 -2675 -1808
rect -2758 -1811 -2601 -1809
rect -2758 -1813 -2752 -1811
rect -2917 -1817 -2752 -1813
rect -2917 -1853 -2913 -1817
rect -2924 -1857 -2899 -1853
rect -2843 -1857 -2839 -1817
rect -2791 -1909 -2786 -1879
rect -2978 -1913 -2786 -1909
rect -3297 -1932 -3176 -1927
rect -3516 -1954 -3451 -1949
rect -3688 -1969 -3588 -1964
rect -3688 -2086 -3684 -1969
rect -3592 -1971 -3588 -1969
rect -3592 -1975 -3514 -1971
rect -3592 -2011 -3588 -1975
rect -3599 -2015 -3574 -2011
rect -3518 -2015 -3514 -1975
rect -3456 -2012 -3451 -1954
rect -3361 -1960 -3289 -1957
rect -3361 -2086 -3356 -1960
rect -3293 -1962 -3289 -1960
rect -3293 -1966 -3215 -1962
rect -3293 -2002 -3289 -1966
rect -3300 -2006 -3275 -2002
rect -3219 -2006 -3215 -1966
rect -2758 -2086 -2752 -1817
rect -2679 -1813 -2601 -1811
rect -2679 -1849 -2675 -1813
rect -2686 -1853 -2661 -1849
rect -2605 -1853 -2601 -1813
rect -2552 -1850 -2547 -1739
rect -2324 -1887 -2311 -1591
rect -2162 -1716 -1775 -1711
rect -2045 -1795 -1835 -1791
rect -2045 -1798 -2036 -1795
rect -2230 -1802 -2036 -1798
rect -2230 -1838 -2226 -1802
rect -2237 -1842 -2212 -1838
rect -2156 -1842 -2152 -1802
rect -2105 -1887 -2100 -1864
rect -2324 -1895 -2100 -1887
rect -2045 -2086 -2036 -1802
rect -1913 -1831 -1909 -1795
rect -1920 -1835 -1895 -1831
rect -1839 -1835 -1835 -1795
rect -1781 -1832 -1775 -1716
rect -4321 -2091 -2036 -2086
<< labels >>
rlabel pdcontact -2859 -1766 -2855 -1756 1 g2n
rlabel space -1766 -792 -1762 -785 1 or1s3
rlabel metal2 -1859 -1307 -1854 -1303 1 c4
rlabel pdcontact -1866 -1295 -1862 -1285 1 c4
rlabel ndcontact -1866 -1315 -1862 -1310 1 c4
rlabel pdcontact -2228 -1428 -2224 -1418 1 or2c4
rlabel ndcontact -2228 -1448 -2224 -1443 1 or2c4
rlabel polycontact -2416 -1139 -2412 -1135 1 p2p1g0
rlabel pdcontact -2368 -1254 -2364 -1244 1 p3p2p1p0c0
rlabel ndcontact -2368 -1274 -2364 -1269 1 p3p2p1p0c0
rlabel polycontact -2417 -1262 -2413 -1258 1 p2p1p0c0
rlabel pdcontact -2364 -1505 -2360 -1495 1 p3p2g1
rlabel ndcontact -2364 -1525 -2360 -1520 1 p3p2g1
rlabel polycontact -2413 -1513 -2409 -1509 1 p2g1
rlabel space -2068 -1651 -2064 -1644 1 or1p3
rlabel pdcontact -2715 -1431 -2711 -1421 1 or2c3
rlabel ndcontact -2715 -1451 -2711 -1446 1 or2c3
rlabel polycontact -2901 -1295 -2897 -1291 1 p1g0
rlabel pdcontact -2853 -1393 -2849 -1383 1 p2p1p0c0
rlabel ndcontact -2853 -1413 -2849 -1408 1 p2p1p0c0
rlabel polycontact -2902 -1401 -2898 -1397 1 p1p0c0
rlabel polycontact -2743 -1667 -2739 -1663 1 or1p2
rlabel ndcontact -2132 -1759 -2128 -1754 1 g3
rlabel pdcontact -2132 -1739 -2128 -1729 1 g3
rlabel polycontact -2851 -1777 -2847 -1773 1 b2
rlabel metal1 -1706 -787 -1695 -783 1 s3
rlabel ndcontact -1710 -795 -1706 -790 1 s3
rlabel pdcontact -1710 -775 -1706 -765 1 s3
rlabel pdiffusion -1769 -778 -1763 -758 1 orpms3
rlabel polycontact -1726 -787 -1722 -783 1 s3n
rlabel ndcontact -1769 -803 -1763 -798 1 s3n
rlabel pdcontact -1759 -778 -1755 -758 1 s3n
rlabel pdcontact -1817 -801 -1813 -791 1 or1s3
rlabel ndcontact -1817 -821 -1813 -816 1 or1s3
rlabel polycontact -1776 -789 -1772 -785 1 or2s3
rlabel ndcontact -1819 -755 -1815 -750 1 or2s3
rlabel pdcontact -1819 -735 -1815 -725 1 or2s3
rlabel ndiffusion -1877 -761 -1871 -751 1 and1nms3
rlabel ndiffusion -1875 -827 -1869 -817 1 and2nms3
rlabel polycontact -1833 -813 -1829 -809 1 and2ns3
rlabel ndcontact -1865 -827 -1861 -817 1 and2ns3
rlabel pdcontact -1874 -798 -1870 -788 1 and2ns3
rlabel polycontact -1835 -747 -1831 -743 1 and1ns3
rlabel ndcontact -1867 -761 -1863 -751 1 and1ns3
rlabel pdcontact -1876 -732 -1872 -722 1 and1ns3
rlabel polycontact -1884 -743 -1880 -739 1 p3not
rlabel pdcontact -1913 -742 -1909 -732 1 p3not
rlabel ndcontact -1913 -762 -1909 -757 1 p3not
rlabel polycontact -1882 -809 -1878 -805 1 c3not
rlabel pdcontact -1913 -798 -1909 -788 1 c3not
rlabel ndcontact -1913 -818 -1909 -813 1 c3not
rlabel polycontact -1868 -743 -1864 -739 1 c3
rlabel polycontact -1929 -810 -1925 -806 1 c3
rlabel polycontact -1866 -809 -1862 -805 1 p3
rlabel polycontact -1929 -754 -1925 -750 1 p3
rlabel metal1 -2328 -805 -2317 -801 1 s2
rlabel pdcontact -2332 -793 -2328 -783 1 s2
rlabel ndcontact -2332 -813 -2328 -808 1 s2
rlabel polycontact -2348 -805 -2344 -801 1 s2n
rlabel ndcontact -2391 -821 -2385 -816 1 s2n
rlabel pdcontact -2381 -796 -2377 -776 1 s2n
rlabel pdiffusion -2391 -796 -2385 -776 1 orpms2
rlabel polycontact -2388 -807 -2384 -803 1 or1s2
rlabel pdcontact -2439 -819 -2435 -809 1 or1s2
rlabel ndcontact -2439 -839 -2435 -834 1 or1s2
rlabel polycontact -2398 -807 -2394 -803 1 or2s2
rlabel ndcontact -2441 -773 -2437 -768 1 or2s2
rlabel pdcontact -2441 -753 -2437 -743 1 or2s2
rlabel polycontact -2455 -831 -2451 -827 1 and2ns2
rlabel ndiffusion -2497 -845 -2491 -835 1 and2nms2
rlabel ndcontact -2487 -845 -2483 -835 1 and2ns2
rlabel pdcontact -2496 -816 -2492 -806 1 and2ns2
rlabel polycontact -2457 -765 -2453 -761 1 and1ns2
rlabel ndcontact -2489 -779 -2485 -769 1 and1ns2
rlabel ndiffusion -2499 -779 -2493 -769 1 and1nms2
rlabel pdcontact -2498 -750 -2494 -740 1 and1ns2
rlabel polycontact -2506 -761 -2502 -757 1 p2not
rlabel pdcontact -2535 -760 -2531 -750 1 p2not
rlabel ndcontact -2535 -780 -2531 -775 1 p2not
rlabel polycontact -2490 -761 -2486 -757 1 c2
rlabel polycontact -2551 -772 -2547 -768 1 p2
rlabel polycontact -2488 -827 -2484 -823 1 p2
rlabel polycontact -2504 -827 -2500 -823 1 c2not
rlabel pdcontact -2535 -816 -2531 -806 1 c2not
rlabel ndcontact -2535 -836 -2531 -831 1 c2not
rlabel polycontact -2551 -828 -2547 -824 1 c2
rlabel pdcontact -2381 -1377 -2377 -1367 1 vdd
rlabel polycontact -2735 -1341 -2731 -1337 1 orc3n
rlabel metal1 -2761 -1349 -2751 -1345 1 orc3n
rlabel ndcontact -2778 -1357 -2772 -1352 1 orc3n
rlabel pdcontact -2768 -1332 -2764 -1312 1 orc3n
rlabel pdcontact -2764 -1434 -2760 -1414 1 or2c3n
rlabel ndcontact -2774 -1459 -2768 -1454 1 or2c3n
rlabel metal1 -2760 -1451 -2751 -1447 1 or2c3n
rlabel polycontact -2731 -1443 -2727 -1439 1 or2c3n
rlabel metal2 -2709 -1443 -2700 -1439 1 or2c3
rlabel polycontact -2659 -1382 -2655 -1378 1 or2c3
rlabel polycontact -2669 -1382 -2665 -1378 1 orc3
rlabel metal1 -2712 -1341 -2702 -1337 1 orc3
rlabel ndcontact -2719 -1349 -2715 -1344 1 orc3
rlabel pdcontact -2719 -1329 -2715 -1319 1 orc3
rlabel ndcontact -1884 -1315 -1880 -1310 1 gnd
rlabel ndcontact -1915 -1323 -1911 -1318 1 gnd
rlabel ndcontact -1933 -1323 -1929 -1318 1 gnd
rlabel pdcontact -1884 -1295 -1880 -1285 1 vdd
rlabel pdcontact -1933 -1298 -1929 -1278 1 vdd
rlabel polycontact -1882 -1307 -1878 -1303 1 coutn
rlabel metal1 -1910 -1315 -1905 -1311 1 coutn
rlabel ndcontact -1925 -1323 -1919 -1318 1 coutn
rlabel pdcontact -1915 -1298 -1911 -1278 1 coutn
rlabel pdiffusion -1925 -1298 -1919 -1278 1 or0pmc4
rlabel polycontact -1932 -1309 -1928 -1305 1 or1c4
rlabel metal1 -2041 -1316 -2033 -1312 1 or1c4
rlabel ndcontact -2051 -1324 -2047 -1319 1 or1c4
rlabel pdcontact -2051 -1304 -2047 -1294 1 or1c4
rlabel polycontact -2067 -1316 -2063 -1312 1 or1c4n
rlabel metal1 -2089 -1324 -2085 -1320 1 or1c4n
rlabel ndcontact -2110 -1332 -2104 -1327 1 or1c4n
rlabel pdcontact -2100 -1307 -2096 -1287 1 or1c4n
rlabel ndcontact -2069 -1324 -2065 -1319 1 gnd
rlabel ndcontact -2100 -1332 -2096 -1327 1 gnd
rlabel ndcontact -2118 -1332 -2114 -1327 1 gnd
rlabel pdcontact -2069 -1304 -2065 -1294 1 vdd
rlabel pdcontact -2118 -1307 -2114 -1287 1 vdd
rlabel pdiffusion -2110 -1307 -2104 -1287 1 or1pmc4
rlabel polycontact -2107 -1318 -2103 -1314 1 or2c4
rlabel metal2 -2204 -1440 -2196 -1436 1 or2c4
rlabel polycontact -2244 -1440 -2240 -1436 1 or2c4n
rlabel metal1 -2270 -1448 -2264 -1444 1 or2c4n
rlabel ndcontact -2287 -1456 -2281 -1451 1 or2c4n
rlabel pdcontact -2277 -1431 -2273 -1411 1 or2c4n
rlabel pdiffusion -2287 -1431 -2281 -1411 1 or2pmc4
rlabel ndcontact -2246 -1448 -2242 -1443 1 gnd
rlabel ndcontact -2277 -1456 -2273 -1451 1 gnd
rlabel ndcontact -2295 -1456 -2291 -1451 1 gnd
rlabel pdcontact -2246 -1428 -2242 -1418 1 vdd
rlabel pdcontact -2295 -1431 -2291 -1411 1 vdd
rlabel polycontact -2117 -1318 -2113 -1314 1 or3c4
rlabel metal1 -2218 -1196 -2213 -1192 1 or3c4
rlabel ndcontact -2227 -1204 -2223 -1199 1 or3c4
rlabel pdcontact -2227 -1184 -2223 -1174 1 or3c4
rlabel polycontact -2243 -1196 -2239 -1192 1 or3nc4
rlabel metal1 -2263 -1204 -2259 -1196 1 or3nc4
rlabel ndcontact -2286 -1212 -2280 -1207 1 or3nc4
rlabel pdcontact -2276 -1187 -2272 -1167 1 or3nc4
rlabel pdiffusion -2286 -1187 -2280 -1167 1 or3pmc4
rlabel ndcontact -2245 -1204 -2241 -1199 1 gnd
rlabel ndcontact -2276 -1212 -2272 -1207 1 gnd
rlabel ndcontact -2294 -1212 -2290 -1207 1 gnd
rlabel pdcontact -2245 -1184 -2241 -1174 1 vdd
rlabel pdcontact -2294 -1187 -2290 -1167 1 vdd
rlabel polycontact -2293 -1198 -2289 -1194 1 p3p2p1g0
rlabel ndcontact -2381 -1397 -2377 -1392 1 gnd
rlabel pdcontact -2382 -1505 -2378 -1495 1 vdd
rlabel ndcontact -2382 -1525 -2378 -1520 1 gnd
rlabel ndcontact -2430 -1531 -2426 -1521 1 gnd
rlabel pdcontact -2412 -1502 -2408 -1492 1 vdd
rlabel pdcontact -2430 -1502 -2426 -1492 1 vdd
rlabel polycontact -2432 -1140 -2428 -1135 1 p3
rlabel metal1 -2354 -1143 -2344 -1139 1 p3p2p1g0
rlabel pdcontact -2367 -1131 -2363 -1121 1 p3p2p1g0
rlabel ndcontact -2367 -1151 -2363 -1146 1 p3p2p1g0
rlabel ndcontact -2385 -1151 -2381 -1146 1 gnd
rlabel ndiffusion -2425 -1157 -2419 -1147 1 and4nmc4
rlabel polycontact -2383 -1143 -2379 -1139 1 p3p2p1g0n
rlabel metal1 -2409 -1147 -2399 -1143 1 p3p2p1g0n
rlabel ndcontact -2415 -1157 -2411 -1147 1 p3p2p1g0n
rlabel pdcontact -2424 -1128 -2420 -1118 1 p3p2p1g0n
rlabel pdcontact -2385 -1131 -2381 -1121 1 vdd
rlabel pdcontact -2415 -1128 -2411 -1118 1 vdd
rlabel pdcontact -2433 -1128 -2429 -1118 1 vdd
rlabel ndcontact -2433 -1157 -2429 -1147 1 gnd
rlabel ndcontact -2434 -1280 -2430 -1270 1 gnd
rlabel ndcontact -2386 -1274 -2382 -1269 1 gnd
rlabel polycontact -2283 -1198 -2279 -1194 1 p3p2p1p0c0
rlabel metal2 -2358 -1266 -2347 -1263 1 p3p2p1p0c0
rlabel polycontact -2384 -1266 -2380 -1262 1 p3p2p1p0c0n
rlabel ndiffusion -2426 -1280 -2420 -1270 1 and3nmc4
rlabel ndcontact -2416 -1280 -2412 -1270 1 p3p2p1p0c0n
rlabel pdcontact -2425 -1251 -2421 -1241 1 p3p2p1p0c0n
rlabel pdcontact -2416 -1251 -2412 -1241 1 vdd
rlabel pdcontact -2434 -1251 -2430 -1241 1 vdd
rlabel pdcontact -2386 -1254 -2382 -1244 1 vdd
rlabel polycontact -2294 -1442 -2290 -1438 1 p3g2
rlabel metal1 -2350 -1389 -2343 -1385 1 p3g2
rlabel ndcontact -2363 -1397 -2359 -1392 1 p3g2
rlabel pdcontact -2363 -1377 -2359 -1367 1 p3g2
rlabel polycontact -2379 -1389 -2375 -1385 1 p3g2n
rlabel metal1 -2403 -1393 -2395 -1389 1 p3g2n
rlabel ndcontact -2411 -1403 -2407 -1393 1 p3g2n
rlabel pdcontact -2420 -1374 -2416 -1364 1 p3g2n
rlabel pdcontact -2411 -1374 -2407 -1364 1 vdd
rlabel pdcontact -2429 -1374 -2425 -1364 1 vdd
rlabel ndcontact -2429 -1403 -2425 -1393 1 gnd
rlabel ndiffusion -2421 -1403 -2415 -1393 1 and2nmc4
rlabel ndiffusion -2422 -1531 -2416 -1521 1 and1nmc4
rlabel metal2 -2352 -1517 -2343 -1514 1 p2p3g1
rlabel polycontact -2380 -1517 -2376 -1513 1 p2p3g1n
rlabel ndcontact -2412 -1531 -2408 -1521 1 p2p3g1n
rlabel pdcontact -2421 -1502 -2417 -1492 1 p2p3g1n
rlabel polycontact -1922 -1309 -1918 -1305 1 g3
rlabel polycontact -2433 -1262 -2429 -1258 1 p3
rlabel polycontact -2428 -1385 -2424 -1381 1 p3
rlabel polycontact -2429 -1513 -2425 -1509 1 p3
rlabel metal1 -2596 -1380 -2591 -1376 1 c3
rlabel ndcontact -2603 -1388 -2599 -1383 1 c3
rlabel pdcontact -2603 -1368 -2599 -1358 1 c3
rlabel polycontact -2619 -1380 -2615 -1376 1 c3n
rlabel metal1 -2639 -1388 -2635 -1376 1 c3n
rlabel ndcontact -2662 -1396 -2656 -1391 1 c3n
rlabel pdcontact -2652 -1371 -2648 -1351 1 c3n
rlabel pdiffusion -2662 -1371 -2656 -1351 1 or1pmc3
rlabel pdiffusion -2774 -1434 -2768 -1414 1 or2pmc3
rlabel polycontact -2771 -1445 -2767 -1441 1 p2g1
rlabel polycontact -2781 -1445 -2777 -1441 1 g2
rlabel pdiffusion -2778 -1332 -2772 -1312 1 or3pmc3
rlabel polycontact -2785 -1343 -2781 -1339 1 p2p1g0
rlabel polycontact -2775 -1343 -2771 -1339 1 p2p1p0c0
rlabel ndiffusion -2910 -1313 -2904 -1303 1 and3nmc3
rlabel metal1 -2848 -1299 -2836 -1295 1 p2p1g0
rlabel ndcontact -2852 -1307 -2848 -1302 1 p2p1g0
rlabel pdcontact -2852 -1287 -2848 -1277 1 p2p1g0
rlabel polycontact -2868 -1299 -2864 -1295 1 p2p1g0n
rlabel ndcontact -2900 -1313 -2896 -1303 1 p2p1g0n
rlabel pdcontact -2909 -1284 -2905 -1274 1 p2p1g0n
rlabel metal2 -2845 -1502 -2834 -1498 1 p2g1
rlabel polycontact -2865 -1502 -2861 -1498 1 p2g1n
rlabel metal1 -2889 -1506 -2881 -1502 1 p2g1n
rlabel ndcontact -2897 -1516 -2893 -1506 1 p2g1n
rlabel pdcontact -2906 -1487 -2902 -1477 1 p2g1n
rlabel ndiffusion -2907 -1516 -2901 -1506 1 and1nmc3
rlabel ndiffusion -2911 -1419 -2905 -1409 1 and2nmc3
rlabel metal2 -2847 -1406 -2837 -1402 1 p2p1p0c0
rlabel polycontact -2869 -1405 -2865 -1401 1 p2p1p0c0n
rlabel ndcontact -2901 -1419 -2897 -1409 1 p2p1p0c0n
rlabel pdcontact -2910 -1390 -2906 -1380 1 p2p1p0c0n
rlabel polycontact -2917 -1295 -2913 -1291 1 p2
rlabel polycontact -2918 -1401 -2914 -1397 1 p2
rlabel polycontact -2914 -1498 -2910 -1494 1 p2
rlabel metal2 -2125 -1751 -2108 -1747 1 g3
rlabel ndiffusion -2190 -1765 -2184 -1755 1 and1nmg3
rlabel polycontact -2148 -1751 -2144 -1747 1 g3n
rlabel ndcontact -2180 -1765 -2176 -1755 1 g3n
rlabel pdcontact -2189 -1736 -2185 -1726 1 g3n
rlabel polycontact -2197 -1747 -2193 -1743 1 a3
rlabel metal1 -2795 -1781 -2780 -1777 1 g2
rlabel pdcontact -2802 -1769 -2798 -1759 1 g2
rlabel ndcontact -2802 -1789 -2798 -1784 1 g2
rlabel ndiffusion -2860 -1795 -2854 -1785 1 and1nmg2
rlabel polycontact -2818 -1781 -2814 -1777 1 g2n
rlabel ndcontact -2850 -1795 -2846 -1785 1 g2n
rlabel polycontact -2867 -1778 -2863 -1773 1 a2
rlabel ndcontact -2820 -1789 -2816 -1784 1 gnd
rlabel ndcontact -2868 -1795 -2864 -1785 1 gnd
rlabel ndcontact -2198 -1765 -2194 -1755 1 gnd
rlabel ndcontact -2150 -1759 -2146 -1754 1 gnd
rlabel metal1 -2156 -1768 -2122 -1765 1 gnd
rlabel metal1 -2204 -1772 -2170 -1769 1 gnd
rlabel metal1 -2826 -1798 -2792 -1795 1 gnd
rlabel metal1 -2874 -1802 -2840 -1799 1 gnd
rlabel metal1 -2826 -1753 -2792 -1749 1 vdd
rlabel metal1 -2874 -1751 -2840 -1747 1 vdd
rlabel metal1 -2204 -1721 -2170 -1717 1 vdd
rlabel metal1 -2156 -1723 -2122 -1719 1 vdd
rlabel pdcontact -2150 -1739 -2146 -1729 1 vdd
rlabel pdcontact -2180 -1736 -2176 -1726 1 vdd
rlabel pdcontact -2198 -1736 -2194 -1726 1 vdd
rlabel pdcontact -2820 -1769 -2816 -1759 1 vdd
rlabel pdcontact -2850 -1766 -2846 -1756 1 vdd
rlabel pdcontact -2868 -1766 -2864 -1756 1 vdd
rlabel pdcontact -2870 -1287 -2866 -1277 1 vdd
rlabel pdcontact -2900 -1284 -2896 -1274 1 vdd
rlabel pdcontact -2918 -1284 -2914 -1274 1 vdd
rlabel pdcontact -2901 -1390 -2897 -1380 1 vdd
rlabel pdcontact -2919 -1390 -2915 -1380 1 vdd
rlabel pdcontact -2897 -1487 -2893 -1477 1 vdd
rlabel pdcontact -2915 -1487 -2911 -1477 1 vdd
rlabel pdcontact -2867 -1490 -2863 -1480 1 vdd
rlabel pdcontact -2871 -1393 -2867 -1383 1 vdd
rlabel pdcontact -2733 -1431 -2729 -1421 1 vdd
rlabel pdcontact -2737 -1329 -2733 -1319 1 vdd
rlabel pdcontact -2786 -1332 -2782 -1312 1 vdd
rlabel pdcontact -2782 -1434 -2778 -1414 1 vdd
rlabel pdcontact -2670 -1371 -2666 -1351 1 vdd
rlabel pdcontact -2621 -1368 -2617 -1358 1 vdd
rlabel ndcontact -2621 -1388 -2617 -1383 1 gnd
rlabel ndcontact -2652 -1396 -2648 -1391 1 gnd
rlabel ndcontact -2670 -1396 -2666 -1391 1 gnd
rlabel ndcontact -2733 -1451 -2729 -1446 1 gnd
rlabel ndcontact -2737 -1349 -2733 -1344 1 gnd
rlabel ndcontact -2768 -1357 -2764 -1352 1 gnd
rlabel ndcontact -2786 -1357 -2782 -1352 1 gnd
rlabel ndcontact -2764 -1459 -2760 -1454 1 gnd
rlabel ndcontact -2782 -1459 -2778 -1454 1 gnd
rlabel ndcontact -2867 -1510 -2863 -1505 1 gnd
rlabel ndcontact -2871 -1413 -2867 -1408 1 gnd
rlabel ndcontact -2870 -1307 -2866 -1302 1 gnd
rlabel ndcontact -2918 -1313 -2914 -1303 1 gnd
rlabel ndcontact -2919 -1419 -2915 -1409 1 gnd
rlabel ndcontact -2915 -1516 -2911 -1506 1 gnd
rlabel metal1 -2873 -1519 -2839 -1516 1 gnd
rlabel metal1 -2921 -1523 -2887 -1520 1 gnd
rlabel metal1 -2876 -1316 -2842 -1313 1 gnd
rlabel metal1 -2924 -1320 -2890 -1317 1 gnd
rlabel metal1 -2925 -1426 -2891 -1423 1 gnd
rlabel metal1 -2877 -1422 -2843 -1419 1 gnd
rlabel metal1 -2739 -1460 -2705 -1457 1 gnd
rlabel metal1 -2788 -1468 -2754 -1465 1 gnd
rlabel metal1 -2743 -1358 -2709 -1355 1 gnd
rlabel metal1 -2792 -1366 -2758 -1363 1 gnd
rlabel metal1 -2676 -1405 -2642 -1402 1 gnd
rlabel metal1 -2627 -1397 -2593 -1394 1 gnd
rlabel metal1 -2388 -1534 -2354 -1531 1 gnd
rlabel metal1 -2436 -1538 -2402 -1535 1 gnd
rlabel metal1 -2387 -1406 -2353 -1403 1 gnd
rlabel metal1 -2435 -1410 -2401 -1407 1 gnd
rlabel metal1 -2392 -1283 -2358 -1280 1 gnd
rlabel metal1 -2440 -1287 -2406 -1284 1 gnd
rlabel metal1 -2391 -1160 -2357 -1157 1 gnd
rlabel metal1 -2439 -1164 -2405 -1161 1 gnd
rlabel metal1 -2251 -1213 -2217 -1210 1 gnd
rlabel metal1 -2300 -1221 -2266 -1218 1 gnd
rlabel metal1 -2252 -1457 -2218 -1454 1 gnd
rlabel metal1 -2301 -1465 -2267 -1462 1 gnd
rlabel metal1 -2124 -1341 -2090 -1338 1 gnd
rlabel metal1 -2075 -1333 -2041 -1330 1 gnd
rlabel metal1 -1939 -1332 -1905 -1329 1 gnd
rlabel metal1 -1890 -1324 -1856 -1321 1 gnd
rlabel metal1 -1890 -1279 -1856 -1275 1 vdd
rlabel metal1 -1939 -1270 -1905 -1266 1 vdd
rlabel metal1 -2075 -1288 -2041 -1284 1 vdd
rlabel metal1 -2124 -1279 -2090 -1275 1 vdd
rlabel metal1 -2251 -1168 -2217 -1164 1 vdd
rlabel metal1 -2300 -1159 -2266 -1155 1 vdd
rlabel metal1 -2391 -1115 -2357 -1111 1 vdd
rlabel metal1 -2439 -1113 -2405 -1109 1 vdd
rlabel metal1 -2392 -1238 -2358 -1234 1 vdd
rlabel metal1 -2440 -1236 -2406 -1232 1 vdd
rlabel metal1 -2252 -1412 -2218 -1408 1 vdd
rlabel metal1 -2301 -1403 -2267 -1399 1 vdd
rlabel metal1 -2388 -1489 -2354 -1485 1 vdd
rlabel metal1 -2436 -1487 -2402 -1483 1 vdd
rlabel metal1 -2387 -1361 -2353 -1357 1 vdd
rlabel metal1 -2435 -1359 -2401 -1355 1 vdd
rlabel metal1 -2627 -1352 -2593 -1348 1 vdd
rlabel metal1 -2676 -1343 -2642 -1339 1 vdd
rlabel metal1 -2739 -1415 -2705 -1411 1 vdd
rlabel metal1 -2788 -1406 -2754 -1402 1 vdd
rlabel metal1 -2743 -1313 -2709 -1309 1 vdd
rlabel metal1 -2792 -1304 -2758 -1300 1 vdd
rlabel metal1 -2873 -1474 -2839 -1470 1 vdd
rlabel metal1 -2921 -1472 -2887 -1468 1 vdd
rlabel metal1 -2877 -1377 -2843 -1373 1 vdd
rlabel metal1 -2925 -1375 -2891 -1371 1 vdd
rlabel metal1 -2876 -1271 -2842 -1267 1 vdd
rlabel metal1 -2924 -1269 -2890 -1265 1 vdd
rlabel metal1 -2008 -1646 -1997 -1642 1 p3
rlabel pdcontact -2012 -1634 -2008 -1624 1 p3
rlabel ndcontact -2012 -1654 -2008 -1649 1 p3
rlabel polycontact -2028 -1646 -2024 -1642 1 outnp3
rlabel pdcontact -2061 -1637 -2057 -1617 1 outnp3
rlabel ndcontact -2071 -1662 -2065 -1657 1 outnp3
rlabel pdiffusion -2071 -1637 -2065 -1617 1 orpmp3
rlabel ndcontact -2119 -1680 -2115 -1675 1 or1p3
rlabel pdcontact -2119 -1660 -2115 -1650 1 or1p3
rlabel ndcontact -2121 -1614 -2117 -1609 1 or2p3
rlabel pdcontact -2121 -1594 -2117 -1584 1 or2p3
rlabel polycontact -2168 -1668 -2164 -1664 1 b3
rlabel ndiffusion -2177 -1686 -2171 -1676 1 and2nmp3
rlabel polycontact -2135 -1672 -2131 -1668 1 and2np3
rlabel ndcontact -2167 -1686 -2163 -1676 1 and2np3
rlabel pdcontact -2176 -1657 -2172 -1647 1 and2np3
rlabel ndiffusion -2179 -1620 -2173 -1610 1 and1nmp3
rlabel polycontact -2170 -1602 -2166 -1598 1 a3
rlabel polycontact -2137 -1606 -2133 -1602 1 and1np3
rlabel ndcontact -2169 -1620 -2165 -1610 1 and1np3
rlabel pdcontact -2178 -1591 -2174 -1581 1 and1np3
rlabel polycontact -2184 -1668 -2180 -1664 1 a3not
rlabel pdcontact -2215 -1657 -2211 -1647 1 a3not
rlabel ndcontact -2215 -1677 -2211 -1672 1 a3not
rlabel polycontact -2231 -1669 -2227 -1665 1 a3
rlabel polycontact -2186 -1602 -2182 -1598 1 b3not
rlabel pdcontact -2215 -1601 -2211 -1591 1 b3not
rlabel ndcontact -2215 -1621 -2211 -1616 1 b3not
rlabel polycontact -2231 -1613 -2227 -1609 1 b3
rlabel metal1 -2683 -1665 -2673 -1661 1 p2
rlabel pdcontact -2687 -1653 -2683 -1643 1 p2
rlabel ndcontact -2687 -1673 -2683 -1668 1 p2
rlabel polycontact -2703 -1665 -2699 -1661 1 outnp2
rlabel pdcontact -2736 -1656 -2732 -1636 1 outnp2
rlabel ndcontact -2746 -1681 -2740 -1676 1 outnp2
rlabel pdiffusion -2746 -1656 -2740 -1636 1 orpmp2
rlabel ndcontact -2794 -1699 -2790 -1694 1 or1p2
rlabel pdcontact -2794 -1679 -2790 -1669 1 or1p2
rlabel polycontact -2753 -1667 -2749 -1663 1 or2p2
rlabel ndcontact -2796 -1633 -2792 -1628 1 or2p2
rlabel pdcontact -2796 -1613 -2792 -1603 1 or2p2
rlabel ndiffusion -2854 -1639 -2848 -1629 1 and1nmp2
rlabel polycontact -2845 -1621 -2841 -1617 1 a2
rlabel polycontact -2812 -1625 -2808 -1621 1 and1np2
rlabel ndcontact -2844 -1639 -2840 -1629 1 and1np2
rlabel pdcontact -2853 -1610 -2849 -1600 1 and1np2
rlabel polycontact -2861 -1621 -2857 -1617 1 b2not
rlabel pdcontact -2890 -1620 -2886 -1610 1 b2not
rlabel ndcontact -2890 -1640 -2886 -1635 1 b2not
rlabel polycontact -2906 -1632 -2902 -1627 1 b2
rlabel ndiffusion -2852 -1705 -2846 -1695 1 and2nmp2
rlabel polycontact -2810 -1691 -2806 -1687 1 and2np2
rlabel ndcontact -2842 -1705 -2838 -1695 1 and2np2
rlabel polycontact -2843 -1687 -2839 -1683 1 b2
rlabel pdcontact -2851 -1676 -2847 -1666 1 and2np2
rlabel polycontact -2859 -1687 -2855 -1683 1 a2not
rlabel pdcontact -2890 -1676 -2886 -1666 1 a2not
rlabel ndcontact -2890 -1696 -2886 -1691 1 a2not
rlabel polycontact -2906 -1688 -2902 -1684 1 a2
rlabel ndcontact -1837 -755 -1833 -750 1 gnd
rlabel metal1 -1843 -764 -1809 -761 1 gnd
rlabel metal1 -1889 -834 -1858 -831 1 gnd
rlabel ndcontact -1885 -761 -1881 -751 1 gnd
rlabel ndcontact -1931 -762 -1927 -757 1 gnd
rlabel metal1 -1891 -768 -1857 -765 1 gnd
rlabel metal1 -1937 -771 -1903 -768 1 gnd
rlabel metal1 -1937 -827 -1903 -824 1 gnd
rlabel ndcontact -1931 -818 -1927 -813 1 gnd
rlabel ndcontact -1835 -821 -1831 -816 1 gnd
rlabel ndcontact -1883 -827 -1879 -817 1 gnd
rlabel metal1 -1841 -830 -1807 -827 1 gnd
rlabel metal1 -1734 -804 -1700 -801 1 gnd
rlabel ndcontact -1728 -795 -1724 -790 1 gnd
rlabel ndcontact -1759 -803 -1755 -798 1 gnd
rlabel ndcontact -1777 -803 -1773 -798 1 gnd
rlabel metal1 -1783 -812 -1749 -809 1 gnd
rlabel pdcontact -1728 -775 -1724 -765 1 vdd
rlabel metal1 -1734 -759 -1700 -755 1 vdd
rlabel pdcontact -1777 -778 -1773 -758 1 vdd
rlabel metal1 -1783 -750 -1749 -746 1 vdd
rlabel pdcontact -1835 -801 -1831 -791 1 vdd
rlabel metal1 -1841 -785 -1807 -781 1 vdd
rlabel pdcontact -1865 -798 -1861 -788 1 vdd
rlabel pdcontact -1883 -798 -1879 -788 1 vdd
rlabel metal1 -1889 -783 -1855 -779 1 vdd
rlabel pdcontact -1931 -798 -1927 -788 1 vdd
rlabel metal1 -1937 -782 -1903 -778 1 vdd
rlabel pdcontact -1837 -735 -1833 -725 1 vdd
rlabel metal1 -1843 -719 -1809 -715 5 vdd
rlabel pdcontact -1867 -732 -1863 -722 1 vdd
rlabel pdcontact -1885 -732 -1881 -722 1 vdd
rlabel metal1 -1891 -717 -1857 -713 5 vdd
rlabel pdcontact -1931 -742 -1927 -732 1 vdd
rlabel metal1 -1937 -726 -1903 -722 1 vdd
rlabel ndcontact -2459 -773 -2455 -768 1 gnd
rlabel metal1 -2465 -782 -2431 -779 1 gnd
rlabel metal1 -2511 -852 -2480 -849 1 gnd
rlabel ndcontact -2507 -779 -2503 -769 1 gnd
rlabel ndcontact -2553 -780 -2549 -775 1 gnd
rlabel metal1 -2513 -786 -2479 -783 1 gnd
rlabel metal1 -2559 -789 -2525 -786 1 gnd
rlabel metal1 -2559 -845 -2525 -842 1 gnd
rlabel ndcontact -2553 -836 -2549 -831 1 gnd
rlabel ndcontact -2457 -839 -2453 -834 1 gnd
rlabel ndcontact -2505 -845 -2501 -835 1 gnd
rlabel metal1 -2463 -848 -2429 -845 1 gnd
rlabel metal1 -2356 -822 -2322 -819 1 gnd
rlabel ndcontact -2350 -813 -2346 -808 1 gnd
rlabel ndcontact -2381 -821 -2377 -816 1 gnd
rlabel ndcontact -2399 -821 -2395 -816 1 gnd
rlabel metal1 -2405 -830 -2371 -827 1 gnd
rlabel pdcontact -2350 -793 -2346 -783 1 vdd
rlabel metal1 -2356 -777 -2322 -773 1 vdd
rlabel pdcontact -2399 -796 -2395 -776 1 vdd
rlabel metal1 -2405 -768 -2371 -764 1 vdd
rlabel pdcontact -2457 -819 -2453 -809 1 vdd
rlabel metal1 -2463 -803 -2429 -799 1 vdd
rlabel pdcontact -2487 -816 -2483 -806 1 vdd
rlabel pdcontact -2505 -816 -2501 -806 1 vdd
rlabel metal1 -2511 -801 -2477 -797 1 vdd
rlabel pdcontact -2553 -816 -2549 -806 1 vdd
rlabel metal1 -2559 -800 -2525 -796 1 vdd
rlabel pdcontact -2459 -753 -2455 -743 1 vdd
rlabel metal1 -2465 -737 -2431 -733 5 vdd
rlabel pdcontact -2489 -750 -2485 -740 1 vdd
rlabel pdcontact -2507 -750 -2503 -740 1 vdd
rlabel metal1 -2513 -735 -2479 -731 5 vdd
rlabel pdcontact -2553 -760 -2549 -750 1 vdd
rlabel metal1 -2559 -744 -2525 -740 1 vdd
rlabel ndcontact -2139 -1614 -2135 -1609 1 gnd
rlabel metal1 -2145 -1623 -2111 -1620 1 gnd
rlabel metal1 -2191 -1693 -2160 -1690 1 gnd
rlabel ndcontact -2187 -1620 -2183 -1610 1 gnd
rlabel ndcontact -2233 -1621 -2229 -1616 1 gnd
rlabel metal1 -2193 -1627 -2159 -1624 1 gnd
rlabel metal1 -2239 -1630 -2205 -1627 1 gnd
rlabel metal1 -2239 -1686 -2205 -1683 1 gnd
rlabel ndcontact -2233 -1677 -2229 -1672 1 gnd
rlabel ndcontact -2137 -1680 -2133 -1675 1 gnd
rlabel ndcontact -2185 -1686 -2181 -1676 1 gnd
rlabel metal1 -2143 -1689 -2109 -1686 1 gnd
rlabel metal1 -2036 -1663 -2002 -1660 1 gnd
rlabel ndcontact -2030 -1654 -2026 -1649 1 gnd
rlabel ndcontact -2061 -1662 -2057 -1657 1 gnd
rlabel ndcontact -2079 -1662 -2075 -1657 1 gnd
rlabel metal1 -2085 -1671 -2051 -1668 1 gnd
rlabel pdcontact -2030 -1634 -2026 -1624 1 vdd
rlabel metal1 -2036 -1618 -2002 -1614 1 vdd
rlabel pdcontact -2079 -1637 -2075 -1617 1 vdd
rlabel metal1 -2085 -1609 -2051 -1605 1 vdd
rlabel pdcontact -2137 -1660 -2133 -1650 1 vdd
rlabel metal1 -2143 -1644 -2109 -1640 1 vdd
rlabel pdcontact -2167 -1657 -2163 -1647 1 vdd
rlabel pdcontact -2185 -1657 -2181 -1647 1 vdd
rlabel metal1 -2191 -1642 -2157 -1638 1 vdd
rlabel pdcontact -2233 -1657 -2229 -1647 1 vdd
rlabel metal1 -2239 -1641 -2205 -1637 1 vdd
rlabel pdcontact -2139 -1594 -2135 -1584 1 vdd
rlabel metal1 -2145 -1578 -2111 -1574 5 vdd
rlabel pdcontact -2169 -1591 -2165 -1581 1 vdd
rlabel pdcontact -2187 -1591 -2183 -1581 1 vdd
rlabel metal1 -2193 -1576 -2159 -1572 5 vdd
rlabel pdcontact -2233 -1601 -2229 -1591 1 vdd
rlabel metal1 -2239 -1585 -2205 -1581 1 vdd
rlabel ndcontact -2814 -1633 -2810 -1628 1 gnd
rlabel metal1 -2820 -1642 -2786 -1639 1 gnd
rlabel metal1 -2866 -1712 -2835 -1709 1 gnd
rlabel ndcontact -2862 -1639 -2858 -1629 1 gnd
rlabel ndcontact -2908 -1640 -2904 -1635 1 gnd
rlabel metal1 -2868 -1646 -2834 -1643 1 gnd
rlabel metal1 -2914 -1649 -2880 -1646 1 gnd
rlabel metal1 -2914 -1705 -2880 -1702 1 gnd
rlabel ndcontact -2908 -1696 -2904 -1691 1 gnd
rlabel ndcontact -2812 -1699 -2808 -1694 1 gnd
rlabel ndcontact -2860 -1705 -2856 -1695 1 gnd
rlabel metal1 -2818 -1708 -2784 -1705 1 gnd
rlabel metal1 -2711 -1682 -2677 -1679 1 gnd
rlabel ndcontact -2705 -1673 -2701 -1668 1 gnd
rlabel ndcontact -2736 -1681 -2732 -1676 1 gnd
rlabel ndcontact -2754 -1681 -2750 -1676 1 gnd
rlabel metal1 -2760 -1690 -2726 -1687 1 gnd
rlabel pdcontact -2705 -1653 -2701 -1643 1 vdd
rlabel metal1 -2711 -1637 -2677 -1633 1 vdd
rlabel pdcontact -2754 -1656 -2750 -1636 1 vdd
rlabel metal1 -2760 -1628 -2726 -1624 1 vdd
rlabel pdcontact -2812 -1679 -2808 -1669 1 vdd
rlabel metal1 -2818 -1663 -2784 -1659 1 vdd
rlabel pdcontact -2842 -1676 -2838 -1666 1 vdd
rlabel pdcontact -2860 -1676 -2856 -1666 1 vdd
rlabel metal1 -2866 -1661 -2832 -1657 1 vdd
rlabel pdcontact -2908 -1676 -2904 -1666 1 vdd
rlabel metal1 -2914 -1660 -2880 -1656 1 vdd
rlabel pdcontact -2814 -1613 -2810 -1603 1 vdd
rlabel metal1 -2820 -1597 -2786 -1593 5 vdd
rlabel pdcontact -2844 -1610 -2840 -1600 1 vdd
rlabel pdcontact -2862 -1610 -2858 -1600 1 vdd
rlabel metal1 -2868 -1595 -2834 -1591 5 vdd
rlabel pdcontact -2908 -1620 -2904 -1610 1 vdd
rlabel metal1 -2914 -1604 -2880 -1600 1 vdd
rlabel polycontact -3363 -1486 -3359 -1482 1 p1g0
rlabel polycontact -3788 -1798 -3784 -1794 1 b0
rlabel polycontact -3211 -787 -3207 -783 1 p1
rlabel polycontact -3817 -1044 -3813 -1040 1 c0
rlabel polycontact -3754 -1099 -3750 -1095 1 c0
rlabel polycontact -3440 -1416 -3436 -1412 1 p1g0n
rlabel pdcontact -3424 -1404 -3420 -1394 1 p1g0
rlabel ndcontact -3424 -1424 -3420 -1419 1 p1g0
rlabel polycontact -3468 -1521 -3464 -1517 1 p1
rlabel polycontact -3473 -1412 -3469 -1408 1 p1
rlabel metal1 -3049 -831 -3038 -827 1 s1
rlabel ndcontact -3053 -839 -3049 -834 1 s1
rlabel pdcontact -3053 -819 -3049 -809 1 s1
rlabel polycontact -3069 -831 -3065 -827 1 s1n
rlabel ndcontact -3112 -847 -3106 -842 1 s1n
rlabel pdcontact -3102 -822 -3098 -802 1 s1n
rlabel pdiffusion -3112 -822 -3106 -802 1 orpms1
rlabel pdcontact -3162 -779 -3158 -769 1 or2s1
rlabel ndcontact -3162 -799 -3158 -794 1 or2s1
rlabel polycontact -3109 -833 -3105 -829 1 or1s1
rlabel polycontact -3119 -833 -3115 -829 1 or2s1
rlabel ndcontact -3160 -865 -3156 -860 1 or1s1
rlabel pdcontact -3160 -845 -3156 -835 1 or1s1
rlabel ndiffusion -3218 -871 -3212 -861 1 and2nms1
rlabel ndiffusion -3220 -805 -3214 -795 1 and1nms1
rlabel polycontact -3178 -791 -3174 -787 1 and1ns1
rlabel polycontact -3176 -857 -3172 -853 1 and2ns1
rlabel ndcontact -3208 -871 -3204 -861 1 and2ns1
rlabel ndcontact -3210 -805 -3206 -795 1 and1ns1
rlabel pdcontact -3219 -776 -3215 -766 1 and1ns1
rlabel pdcontact -3217 -842 -3213 -832 1 and2ns1
rlabel polycontact -3209 -853 -3205 -849 1 c1
rlabel polycontact -3225 -853 -3221 -849 1 p1not
rlabel pdcontact -3256 -842 -3252 -832 1 p1not
rlabel ndcontact -3256 -862 -3252 -857 1 p1not
rlabel polycontact -3227 -787 -3223 -783 1 c1not
rlabel pdcontact -3256 -786 -3252 -776 1 c1not
rlabel ndcontact -3256 -806 -3252 -801 1 c1not
rlabel polycontact -3272 -798 -3268 -794 1 c1
rlabel polycontact -3772 -1033 -3768 -1029 1 cinnot
rlabel pdcontact -3801 -1032 -3797 -1022 1 cinnot
rlabel ndcontact -3801 -1052 -3797 -1047 1 cinnot
rlabel polycontact -3272 -854 -3268 -850 1 p1
rlabel metal1 -3594 -1077 -3583 -1073 1 s0
rlabel ndcontact -3598 -1085 -3594 -1080 1 s0
rlabel pdcontact -3598 -1065 -3594 -1055 1 s0
rlabel polycontact -3614 -1077 -3610 -1073 1 s0n
rlabel pdcontact -3647 -1068 -3643 -1048 1 s0n
rlabel ndcontact -3657 -1093 -3651 -1088 1 s0n
rlabel pdiffusion -3657 -1068 -3651 -1048 1 orpms0
rlabel polycontact -3664 -1079 -3660 -1075 1 or2s0
rlabel polycontact -3654 -1079 -3650 -1075 1 or1s0
rlabel pdcontact -3705 -1091 -3701 -1081 1 or1s0
rlabel ndcontact -3705 -1111 -3701 -1106 1 or1s0
rlabel ndcontact -3707 -1045 -3703 -1040 1 or2s0
rlabel pdcontact -3707 -1025 -3703 -1015 1 or2s0
rlabel polycontact -3723 -1037 -3719 -1033 1 and1ns0
rlabel pdcontact -3764 -1022 -3760 -1012 1 and1ns0
rlabel ndcontact -3755 -1051 -3751 -1041 1 and1ns0
rlabel ndiffusion -3765 -1051 -3759 -1041 1 and1nms0
rlabel ndiffusion -3763 -1117 -3757 -1107 1 and2nms0
rlabel polycontact -3721 -1103 -3717 -1099 1 and2ns0
rlabel ndcontact -3753 -1117 -3749 -1107 1 and2ns0
rlabel pdcontact -3762 -1088 -3758 -1078 1 and2ns0
rlabel ndcontact -3801 -1108 -3797 -1103 1 p0not
rlabel pdcontact -3801 -1088 -3797 -1078 1 p0not
rlabel polycontact -3770 -1099 -3766 -1095 1 p0not
rlabel polycontact -3756 -1033 -3752 -1029 1 p0
rlabel polycontact -3817 -1100 -3813 -1096 1 p0
rlabel polycontact -3248 -1476 -3244 -1472 1 or1c2
rlabel metal1 -3286 -1484 -3282 -1472 1 or1c2
rlabel ndcontact -3297 -1492 -3293 -1487 1 or1c2
rlabel pdcontact -3297 -1472 -3293 -1462 1 or1c2
rlabel polycontact -3313 -1484 -3309 -1480 1 or1c2n
rlabel metal1 -3341 -1492 -3329 -1488 1 or1c2n
rlabel ndcontact -3356 -1500 -3350 -1495 1 or1c2n
rlabel pdcontact -3346 -1475 -3342 -1455 1 or1c2n
rlabel polycontact -3484 -1521 -3480 -1517 1 p0c0
rlabel polycontact -3719 -1534 -3715 -1530 1 p0c0
rlabel metal1 -3754 -1534 -3745 -1530 1 p0c0
rlabel ndcontact -3758 -1542 -3754 -1537 1 p0c0
rlabel pdcontact -3758 -1522 -3754 -1512 1 p0c0
rlabel polycontact -3774 -1534 -3770 -1530 1 p0c0n
rlabel metal1 -3800 -1538 -3790 -1534 1 p0c0n
rlabel ndcontact -3806 -1548 -3802 -1538 1 p0c0n
rlabel pdcontact -3815 -1519 -3811 -1509 1 p0c0n
rlabel ndiffusion -3816 -1548 -3810 -1538 1 andnmc1
rlabel ndiffusion -3482 -1430 -3476 -1420 1 and2nmc2
rlabel ndiffusion -3477 -1539 -3471 -1529 1 and1nmc2
rlabel metal1 -3459 -1529 -3451 -1525 1 p1p0c0n
rlabel pdcontact -3476 -1510 -3472 -1500 1 p1p0c0n
rlabel ndcontact -3467 -1539 -3463 -1529 1 p1p0c0n
rlabel polycontact -3435 -1525 -3431 -1521 1 p1p0c0n
rlabel metal1 -3415 -1525 -3406 -1521 1 p1p0c0
rlabel pdcontact -3419 -1513 -3415 -1503 1 p1p0c0
rlabel ndcontact -3419 -1533 -3415 -1528 1 p1p0c0
rlabel polycontact -3353 -1486 -3349 -1482 1 p1p0c0
rlabel metal3 -3424 -1416 -3412 -1412 1 p1g0
rlabel ndcontact -3472 -1430 -3468 -1420 1 p1g0n
rlabel pdcontact -3481 -1401 -3477 -1391 1 p1g0n
rlabel polycontact -3489 -1413 -3485 -1408 1 g0
rlabel pdiffusion -3356 -1475 -3350 -1455 1 or1pmc2
rlabel pdiffusion -3241 -1465 -3235 -1445 1 or2pmc2
rlabel pdcontact -3231 -1465 -3227 -1445 1 c2n
rlabel ndcontact -3241 -1490 -3235 -1485 1 c2n
rlabel polycontact -3198 -1474 -3194 -1470 1 c2n
rlabel metal1 -3168 -1474 -3156 -1470 1 c2
rlabel pdcontact -3182 -1462 -3178 -1452 1 c2
rlabel ndcontact -3182 -1482 -3178 -1477 1 c2
rlabel polycontact -3238 -1476 -3234 -1472 1 g1
rlabel ndcontact -3653 -1540 -3649 -1535 1 c1
rlabel pdcontact -3653 -1520 -3649 -1510 1 c1
rlabel polycontact -3669 -1532 -3665 -1528 1 c1n
rlabel ndcontact -3712 -1548 -3706 -1543 1 c1n
rlabel pdcontact -3702 -1523 -3698 -1503 1 c1n
rlabel pdiffusion -3712 -1523 -3706 -1503 1 orpmc1
rlabel polycontact -3709 -1534 -3705 -1530 1 g0
rlabel polycontact -3823 -1530 -3819 -1526 1 p0
rlabel metal3 -3891 -1475 -3873 -1469 1 c0
rlabel metal1 -3345 -1782 -3328 -1778 1 g1
rlabel ndcontact -3352 -1790 -3348 -1785 1 g1
rlabel pdcontact -3352 -1770 -3348 -1760 1 g1
rlabel polycontact -3368 -1782 -3364 -1778 1 g1n
rlabel ndiffusion -3410 -1796 -3404 -1786 1 and1nmg1
rlabel ndcontact -3400 -1796 -3396 -1786 1 g1n
rlabel pdcontact -3409 -1767 -3405 -1757 1 g1n
rlabel polycontact -3401 -1778 -3397 -1774 1 b1
rlabel polycontact -3417 -1779 -3413 -1774 1 a1
rlabel metal1 -3733 -1803 -3720 -1798 1 g0
rlabel ndcontact -3739 -1810 -3735 -1805 1 g0
rlabel pdcontact -3739 -1790 -3735 -1780 1 g0
rlabel ndiffusion -3797 -1816 -3791 -1806 1 and1nmg0
rlabel ndcontact -3787 -1816 -3783 -1806 1 g0n
rlabel pdcontact -3796 -1787 -3792 -1777 1 g0n
rlabel polycontact -3755 -1802 -3751 -1798 1 g0n
rlabel polycontact -3804 -1799 -3800 -1794 1 a0
rlabel ndcontact -3757 -1810 -3753 -1805 1 gnd
rlabel ndcontact -3805 -1816 -3801 -1806 1 gnd
rlabel ndcontact -3418 -1796 -3414 -1786 1 gnd
rlabel ndcontact -3370 -1790 -3366 -1785 1 gnd
rlabel metal1 -3376 -1799 -3342 -1796 1 gnd
rlabel metal1 -3424 -1803 -3390 -1800 1 gnd
rlabel metal1 -3763 -1819 -3729 -1816 1 gnd
rlabel metal1 -3811 -1823 -3777 -1820 1 gnd
rlabel metal1 -3763 -1774 -3729 -1770 1 vdd
rlabel metal1 -3811 -1772 -3777 -1768 1 vdd
rlabel metal1 -3424 -1752 -3390 -1748 1 vdd
rlabel metal1 -3376 -1754 -3342 -1750 1 vdd
rlabel pdcontact -3370 -1770 -3366 -1760 1 vdd
rlabel pdcontact -3400 -1767 -3396 -1757 1 vdd
rlabel pdcontact -3418 -1767 -3414 -1757 1 vdd
rlabel pdcontact -3757 -1790 -3753 -1780 1 vdd
rlabel pdcontact -3787 -1787 -3783 -1777 1 vdd
rlabel pdcontact -3805 -1787 -3801 -1777 1 vdd
rlabel pdcontact -3249 -1465 -3245 -1445 1 vdd
rlabel pdcontact -3364 -1475 -3360 -1455 1 vdd
rlabel pdcontact -3720 -1523 -3716 -1503 1 vdd
rlabel pdcontact -3671 -1520 -3667 -1510 1 vdd
rlabel pdcontact -3776 -1522 -3772 -1512 1 vdd
rlabel pdcontact -3806 -1519 -3802 -1509 1 vdd
rlabel pdcontact -3824 -1519 -3820 -1509 1 vdd
rlabel pdcontact -3442 -1404 -3438 -1394 1 vdd
rlabel pdcontact -3472 -1401 -3468 -1391 1 vdd
rlabel pdcontact -3490 -1401 -3486 -1391 1 vdd
rlabel pdcontact -3467 -1510 -3463 -1500 1 vdd
rlabel pdcontact -3485 -1510 -3481 -1500 1 vdd
rlabel pdcontact -3437 -1513 -3433 -1503 1 vdd
rlabel pdcontact -3315 -1472 -3311 -1462 1 vdd
rlabel pdcontact -3200 -1462 -3196 -1452 1 vdd
rlabel ndcontact -3200 -1482 -3196 -1477 1 gnd
rlabel ndcontact -3231 -1490 -3227 -1485 1 gnd
rlabel ndcontact -3249 -1490 -3245 -1485 1 gnd
rlabel ndcontact -3315 -1492 -3311 -1487 1 gnd
rlabel ndcontact -3346 -1500 -3342 -1495 1 gnd
rlabel ndcontact -3364 -1500 -3360 -1495 1 gnd
rlabel ndcontact -3437 -1533 -3433 -1528 1 gnd
rlabel ndcontact -3442 -1424 -3438 -1419 1 gnd
rlabel ndcontact -3490 -1430 -3486 -1420 1 gnd
rlabel ndcontact -3485 -1539 -3481 -1529 1 gnd
rlabel ndcontact -3671 -1540 -3667 -1535 1 gnd
rlabel ndcontact -3702 -1548 -3698 -1543 1 gnd
rlabel ndcontact -3720 -1548 -3716 -1543 1 gnd
rlabel ndcontact -3776 -1542 -3772 -1537 1 gnd
rlabel ndcontact -3824 -1548 -3820 -1538 1 gnd
rlabel metal1 -3830 -1555 -3796 -1552 1 gnd
rlabel metal1 -3782 -1551 -3748 -1548 1 gnd
rlabel metal1 -3726 -1557 -3692 -1554 1 gnd
rlabel metal1 -3677 -1549 -3643 -1546 1 gnd
rlabel metal1 -3448 -1433 -3414 -1430 1 gnd
rlabel metal1 -3496 -1437 -3462 -1434 1 gnd
rlabel metal1 -3491 -1546 -3457 -1543 1 gnd
rlabel metal1 -3443 -1542 -3409 -1539 1 gnd
rlabel metal1 -3370 -1509 -3336 -1506 1 gnd
rlabel metal1 -3321 -1501 -3287 -1498 1 gnd
rlabel metal1 -3255 -1499 -3221 -1496 1 gnd
rlabel metal1 -3206 -1491 -3172 -1488 1 gnd
rlabel metal1 -3206 -1446 -3172 -1442 1 vdd
rlabel metal1 -3255 -1437 -3221 -1433 1 vdd
rlabel metal1 -3321 -1456 -3287 -1452 1 vdd
rlabel metal1 -3370 -1447 -3336 -1443 1 vdd
rlabel metal1 -3443 -1497 -3409 -1493 1 vdd
rlabel metal1 -3491 -1495 -3457 -1491 1 vdd
rlabel metal1 -3448 -1388 -3414 -1384 1 vdd
rlabel metal1 -3496 -1386 -3462 -1382 1 vdd
rlabel metal1 -3677 -1504 -3643 -1500 1 vdd
rlabel metal1 -3726 -1495 -3692 -1491 1 vdd
rlabel metal1 -3782 -1506 -3748 -1502 1 vdd
rlabel metal1 -3830 -1504 -3796 -1500 1 vdd
rlabel metal1 -3280 -770 -3246 -766 1 vdd
rlabel pdcontact -3274 -786 -3270 -776 1 vdd
rlabel metal1 -3234 -761 -3200 -757 5 vdd
rlabel pdcontact -3228 -776 -3224 -766 1 vdd
rlabel pdcontact -3210 -776 -3206 -766 1 vdd
rlabel metal1 -3186 -763 -3152 -759 5 vdd
rlabel pdcontact -3180 -779 -3176 -769 1 vdd
rlabel metal1 -3280 -826 -3246 -822 1 vdd
rlabel pdcontact -3274 -842 -3270 -832 1 vdd
rlabel metal1 -3232 -827 -3198 -823 1 vdd
rlabel pdcontact -3226 -842 -3222 -832 1 vdd
rlabel pdcontact -3208 -842 -3204 -832 1 vdd
rlabel metal1 -3184 -829 -3150 -825 1 vdd
rlabel pdcontact -3178 -845 -3174 -835 1 vdd
rlabel metal1 -3126 -794 -3092 -790 1 vdd
rlabel pdcontact -3120 -822 -3116 -802 1 vdd
rlabel metal1 -3077 -803 -3043 -799 1 vdd
rlabel pdcontact -3071 -819 -3067 -809 1 vdd
rlabel metal1 -3126 -856 -3092 -853 1 gnd
rlabel ndcontact -3120 -847 -3116 -842 1 gnd
rlabel ndcontact -3102 -847 -3098 -842 1 gnd
rlabel ndcontact -3071 -839 -3067 -834 1 gnd
rlabel metal1 -3077 -848 -3043 -845 1 gnd
rlabel metal1 -3184 -874 -3150 -871 1 gnd
rlabel ndcontact -3226 -871 -3222 -861 1 gnd
rlabel ndcontact -3178 -865 -3174 -860 1 gnd
rlabel ndcontact -3274 -862 -3270 -857 1 gnd
rlabel metal1 -3280 -871 -3246 -868 1 gnd
rlabel metal1 -3280 -815 -3246 -812 1 gnd
rlabel metal1 -3234 -812 -3200 -809 1 gnd
rlabel ndcontact -3274 -806 -3270 -801 1 gnd
rlabel ndcontact -3228 -805 -3224 -795 1 gnd
rlabel metal1 -3232 -878 -3201 -875 1 gnd
rlabel metal1 -3186 -808 -3152 -805 1 gnd
rlabel ndcontact -3180 -799 -3176 -794 1 gnd
rlabel ndcontact -3725 -1045 -3721 -1040 1 gnd
rlabel metal1 -3731 -1054 -3697 -1051 1 gnd
rlabel metal1 -3777 -1124 -3746 -1121 1 gnd
rlabel ndcontact -3773 -1051 -3769 -1041 1 gnd
rlabel ndcontact -3819 -1052 -3815 -1047 1 gnd
rlabel metal1 -3779 -1058 -3745 -1055 1 gnd
rlabel metal1 -3825 -1061 -3791 -1058 1 gnd
rlabel metal1 -3825 -1117 -3791 -1114 1 gnd
rlabel ndcontact -3819 -1108 -3815 -1103 1 gnd
rlabel ndcontact -3723 -1111 -3719 -1106 1 gnd
rlabel ndcontact -3771 -1117 -3767 -1107 1 gnd
rlabel metal1 -3729 -1120 -3695 -1117 1 gnd
rlabel metal1 -3622 -1094 -3588 -1091 1 gnd
rlabel ndcontact -3616 -1085 -3612 -1080 1 gnd
rlabel ndcontact -3647 -1093 -3643 -1088 1 gnd
rlabel ndcontact -3665 -1093 -3661 -1088 1 gnd
rlabel metal1 -3671 -1102 -3637 -1099 1 gnd
rlabel pdcontact -3616 -1065 -3612 -1055 1 vdd
rlabel metal1 -3622 -1049 -3588 -1045 1 vdd
rlabel pdcontact -3665 -1068 -3661 -1048 1 vdd
rlabel metal1 -3671 -1040 -3637 -1036 1 vdd
rlabel pdcontact -3723 -1091 -3719 -1081 1 vdd
rlabel metal1 -3729 -1075 -3695 -1071 1 vdd
rlabel pdcontact -3753 -1088 -3749 -1078 1 vdd
rlabel pdcontact -3771 -1088 -3767 -1078 1 vdd
rlabel metal1 -3777 -1073 -3743 -1069 1 vdd
rlabel pdcontact -3819 -1088 -3815 -1078 1 vdd
rlabel metal1 -3825 -1072 -3791 -1068 1 vdd
rlabel pdcontact -3725 -1025 -3721 -1015 1 vdd
rlabel metal1 -3731 -1009 -3697 -1005 5 vdd
rlabel pdcontact -3755 -1022 -3751 -1012 1 vdd
rlabel pdcontact -3773 -1022 -3769 -1012 1 vdd
rlabel metal1 -3779 -1007 -3745 -1003 5 vdd
rlabel pdcontact -3819 -1032 -3815 -1022 1 vdd
rlabel metal1 -3825 -1016 -3791 -1012 1 vdd
rlabel metal1 -3244 -1665 -3233 -1661 1 p1
rlabel ndcontact -3248 -1673 -3244 -1668 1 p1
rlabel pdcontact -3248 -1653 -3244 -1643 1 p1
rlabel polycontact -3264 -1665 -3260 -1661 1 outnp1
rlabel ndcontact -3307 -1681 -3301 -1676 1 outnp1
rlabel pdcontact -3297 -1656 -3293 -1636 1 outnp1
rlabel pdiffusion -3307 -1656 -3301 -1636 1 orpmp1
rlabel pdcontact -3357 -1613 -3353 -1603 1 or2p1
rlabel ndcontact -3357 -1633 -3353 -1628 1 or2p1
rlabel polycontact -3314 -1667 -3310 -1663 1 or2p1
rlabel polycontact -3304 -1667 -3300 -1663 1 or1p1
rlabel pdcontact -3355 -1679 -3351 -1669 1 or1p1
rlabel ndcontact -3355 -1699 -3351 -1694 1 or1p1
rlabel polycontact -3371 -1691 -3367 -1687 1 and2np1
rlabel ndiffusion -3413 -1705 -3407 -1695 1 and2nmp1
rlabel ndcontact -3403 -1705 -3399 -1695 1 and2np1
rlabel pdcontact -3412 -1676 -3408 -1666 1 and2np1
rlabel polycontact -3404 -1687 -3400 -1683 1 b1
rlabel polycontact -3406 -1621 -3402 -1617 1 a1
rlabel polycontact -3373 -1625 -3369 -1621 1 and1np1
rlabel ndiffusion -3415 -1639 -3409 -1629 1 and1nmp1
rlabel ndcontact -3405 -1639 -3401 -1629 1 and1np1
rlabel pdcontact -3414 -1610 -3410 -1600 1 and1np1
rlabel pdcontact -3451 -1620 -3447 -1610 1 b1not
rlabel ndcontact -3451 -1640 -3447 -1635 1 b1not
rlabel polycontact -3422 -1621 -3418 -1617 1 b1not
rlabel polycontact -3420 -1687 -3416 -1683 1 a1not
rlabel pdcontact -3451 -1676 -3447 -1666 1 a1not
rlabel ndcontact -3451 -1696 -3447 -1691 1 a1not
rlabel polycontact -3467 -1688 -3463 -1684 1 a1
rlabel polycontact -3467 -1632 -3463 -1628 1 b1
rlabel pdcontact -3600 -1655 -3596 -1645 1 p0
rlabel ndcontact -3600 -1675 -3596 -1670 1 p0
rlabel polycontact -3616 -1667 -3612 -1663 1 outnp0
rlabel ndcontact -3659 -1683 -3653 -1678 1 outnp0
rlabel pdcontact -3649 -1658 -3645 -1638 1 outnp0
rlabel pdiffusion -3659 -1658 -3653 -1638 1 orpmp0
rlabel polycontact -3656 -1669 -3652 -1665 1 or1p0
rlabel polycontact -3666 -1669 -3662 -1665 1 or2p0
rlabel ndcontact -3709 -1635 -3705 -1630 1 or2p0
rlabel pdcontact -3709 -1615 -3705 -1605 1 or2p0
rlabel pdcontact -3707 -1681 -3703 -1671 1 or1p0
rlabel ndcontact -3707 -1701 -3703 -1696 1 or1p0
rlabel polycontact -3723 -1693 -3719 -1689 1 and2np0
rlabel polycontact -3725 -1627 -3721 -1623 1 and1np0
rlabel pdcontact -3766 -1612 -3762 -1602 1 and1np0
rlabel ndiffusion -3767 -1641 -3761 -1631 1 and1nmp0
rlabel ndcontact -3757 -1641 -3753 -1631 1 and1np0
rlabel ndcontact -3755 -1707 -3751 -1697 1 and2np0
rlabel pdcontact -3764 -1678 -3760 -1668 1 and2np0
rlabel ndiffusion -3765 -1707 -3759 -1697 1 and2nmp0
rlabel metal1 -3596 -1667 -3585 -1663 1 p0
rlabel polycontact -3756 -1689 -3752 -1685 1 b0
rlabel polycontact -3758 -1623 -3754 -1619 1 a0
rlabel polycontact -3774 -1623 -3770 -1619 1 b0not
rlabel polycontact -3772 -1689 -3768 -1685 1 a0not
rlabel ndcontact -3803 -1642 -3799 -1637 1 b0not
rlabel ndcontact -3803 -1698 -3799 -1693 1 a0not
rlabel polycontact -3819 -1690 -3815 -1686 1 a0
rlabel polycontact -3819 -1634 -3815 -1630 1 b0
rlabel ndcontact -3727 -1635 -3723 -1630 1 gnd
rlabel metal1 -3733 -1644 -3699 -1641 1 gnd
rlabel metal1 -3779 -1714 -3748 -1711 1 gnd
rlabel pdcontact -3803 -1678 -3799 -1668 1 anot
rlabel pdcontact -3803 -1622 -3799 -1612 1 bnot
rlabel ndcontact -3775 -1641 -3771 -1631 1 gnd
rlabel ndcontact -3821 -1642 -3817 -1637 1 gnd
rlabel metal1 -3781 -1648 -3747 -1645 1 gnd
rlabel metal1 -3827 -1651 -3793 -1648 1 gnd
rlabel metal1 -3827 -1707 -3793 -1704 1 gnd
rlabel ndcontact -3821 -1698 -3817 -1693 1 gnd
rlabel ndcontact -3725 -1701 -3721 -1696 1 gnd
rlabel ndcontact -3773 -1707 -3769 -1697 1 gnd
rlabel metal1 -3731 -1710 -3697 -1707 1 gnd
rlabel metal1 -3624 -1684 -3590 -1681 1 gnd
rlabel ndcontact -3618 -1675 -3614 -1670 1 gnd
rlabel ndcontact -3649 -1683 -3645 -1678 1 gnd
rlabel ndcontact -3667 -1683 -3663 -1678 1 gnd
rlabel metal1 -3673 -1692 -3639 -1689 1 gnd
rlabel pdcontact -3618 -1655 -3614 -1645 1 vdd
rlabel metal1 -3624 -1639 -3590 -1635 1 vdd
rlabel pdcontact -3667 -1658 -3663 -1638 1 vdd
rlabel metal1 -3673 -1630 -3639 -1626 1 vdd
rlabel pdcontact -3725 -1681 -3721 -1671 1 vdd
rlabel metal1 -3731 -1665 -3697 -1661 1 vdd
rlabel pdcontact -3755 -1678 -3751 -1668 1 vdd
rlabel pdcontact -3773 -1678 -3769 -1668 1 vdd
rlabel metal1 -3779 -1663 -3745 -1659 1 vdd
rlabel pdcontact -3821 -1678 -3817 -1668 1 vdd
rlabel metal1 -3827 -1662 -3793 -1658 1 vdd
rlabel pdcontact -3727 -1615 -3723 -1605 1 vdd
rlabel metal1 -3733 -1599 -3699 -1595 5 vdd
rlabel pdcontact -3757 -1612 -3753 -1602 1 vdd
rlabel pdcontact -3775 -1612 -3771 -1602 1 vdd
rlabel metal1 -3781 -1597 -3747 -1593 5 vdd
rlabel pdcontact -3821 -1622 -3817 -1612 1 vdd
rlabel metal1 -3827 -1606 -3793 -1602 1 vdd
rlabel ndcontact -3375 -1633 -3371 -1628 1 gnd
rlabel metal1 -3381 -1642 -3347 -1639 1 gnd
rlabel metal1 -3427 -1712 -3396 -1709 1 gnd
rlabel ndcontact -3423 -1639 -3419 -1629 1 gnd
rlabel ndcontact -3469 -1640 -3465 -1635 1 gnd
rlabel metal1 -3429 -1646 -3395 -1643 1 gnd
rlabel metal1 -3475 -1649 -3441 -1646 1 gnd
rlabel metal1 -3475 -1705 -3441 -1702 1 gnd
rlabel ndcontact -3469 -1696 -3465 -1691 1 gnd
rlabel ndcontact -3373 -1699 -3369 -1694 1 gnd
rlabel ndcontact -3421 -1705 -3417 -1695 1 gnd
rlabel metal1 -3379 -1708 -3345 -1705 1 gnd
rlabel metal1 -3272 -1682 -3238 -1679 1 gnd
rlabel ndcontact -3266 -1673 -3262 -1668 1 gnd
rlabel ndcontact -3297 -1681 -3293 -1676 1 gnd
rlabel ndcontact -3315 -1681 -3311 -1676 1 gnd
rlabel metal1 -3321 -1690 -3287 -1687 1 gnd
rlabel pdcontact -3266 -1653 -3262 -1643 1 vdd
rlabel metal1 -3272 -1637 -3238 -1633 1 vdd
rlabel pdcontact -3315 -1656 -3311 -1636 1 vdd
rlabel metal1 -3321 -1628 -3287 -1624 1 vdd
rlabel pdcontact -3373 -1679 -3369 -1669 1 vdd
rlabel metal1 -3379 -1663 -3345 -1659 1 vdd
rlabel pdcontact -3403 -1676 -3399 -1666 1 vdd
rlabel pdcontact -3421 -1676 -3417 -1666 1 vdd
rlabel metal1 -3427 -1661 -3393 -1657 1 vdd
rlabel pdcontact -3469 -1676 -3465 -1666 1 vdd
rlabel metal1 -3475 -1660 -3441 -1656 1 vdd
rlabel pdcontact -3375 -1613 -3371 -1603 1 vdd
rlabel metal1 -3381 -1597 -3347 -1593 5 vdd
rlabel pdcontact -3405 -1610 -3401 -1600 1 vdd
rlabel pdcontact -3423 -1610 -3419 -1600 1 vdd
rlabel metal1 -3429 -1595 -3395 -1591 5 vdd
rlabel pdcontact -3469 -1620 -3465 -1610 1 vdd
rlabel metal1 -3475 -1604 -3441 -1600 1 vdd
rlabel metal1 -2050 -1654 -2044 -1650 1 outnp3
rlabel polycontact -2078 -1648 -2074 -1644 1 or2p3
rlabel metal2 -2105 -1651 -2096 -1648 1 or1p3
rlabel metal1 -2117 -1606 -2108 -1602 1 or2p3
rlabel pdcontact -2849 -1490 -2845 -1480 1 p2g1
rlabel ndcontact -2849 -1510 -2845 -1505 1 p2g1
rlabel metal2 -2111 -1672 -2100 -1668 1 or1p3
rlabel metal2 -1806 -813 -1798 -809 1 or1s3
rlabel polycontact -3807 -1530 -3803 -1526 1 c0
rlabel polycontact -2898 -1498 -2894 -1494 1 g1
rlabel polycontact -2412 -1385 -2408 -1381 1 g2
rlabel polysilicon -3705 -1534 -3703 -1530 1 g0
rlabel polysilicon -3234 -1476 -3232 -1472 1 g1
rlabel polysilicon -2900 -1498 -2898 -1494 1 g1
rlabel polysilicon -2414 -1385 -2412 -1381 1 g2
rlabel polysilicon -1918 -1309 -1916 -1305 1 g3
rlabel polysilicon -2064 -1648 -2062 -1644 1 or1p3
rlabel polysilicon -1762 -789 -1760 -785 1 or1s3
rlabel polysilicon -3809 -1530 -3807 -1526 1 c0
rlabel polysilicon -2279 -1198 -2277 -1194 1 p3p2p1p0c0
rlabel polycontact -2284 -1442 -2280 -1438 1 p3p2g1
rlabel polysilicon -2280 -1442 -2278 -1438 1 p3p2g1
rlabel metal1 -4310 -1315 -4278 -1312 5 vdd
rlabel pdcontact -4304 -1339 -4300 -1319 1 vdd
rlabel metal1 -4310 -1371 -4278 -1368 1 gnd
rlabel ndcontact -4304 -1363 -4300 -1358 1 gnd
rlabel polycontact -4280 -1352 -4276 -1348 1 clk
rlabel metal1 -4258 -1315 -4234 -1312 5 vdd
rlabel pdcontact -4252 -1339 -4248 -1329 1 vdd
rlabel metal1 -4263 -1392 -4229 -1387 1 gnd
rlabel ndcontact -4237 -1374 -4233 -1364 1 gnd
rlabel polycontact -4251 -1352 -4247 -1348 1 clk
rlabel metal1 -4224 -1315 -4200 -1312 1 vdd
rlabel pdcontact -4218 -1332 -4214 -1322 1 vdd
rlabel ndcontact -4218 -1374 -4214 -1364 1 gnd
rlabel metal1 -4221 -1390 -4197 -1385 1 gnd
rlabel polycontact -4195 -1356 -4191 -1352 1 clk
rlabel metal1 -4180 -1336 -4146 -1332 1 vdd
rlabel pdcontact -4174 -1352 -4170 -1342 1 vdd
rlabel ndcontact -4174 -1372 -4170 -1367 1 gnd
rlabel metal1 -4180 -1381 -4146 -1378 1 gnd
rlabel metal1 -3857 -567 -3825 -564 5 vdd
rlabel pdcontact -3851 -591 -3847 -571 1 vdd
rlabel metal1 -3857 -623 -3825 -620 1 gnd
rlabel ndcontact -3851 -615 -3847 -610 1 gnd
rlabel polycontact -3827 -604 -3823 -600 1 clk
rlabel metal1 -3805 -567 -3781 -564 5 vdd
rlabel pdcontact -3799 -591 -3795 -581 1 vdd
rlabel metal1 -3810 -644 -3776 -639 1 gnd
rlabel ndcontact -3784 -626 -3780 -616 1 gnd
rlabel polycontact -3798 -604 -3794 -600 1 clk
rlabel metal1 -3771 -567 -3747 -564 1 vdd
rlabel pdcontact -3765 -584 -3761 -574 1 vdd
rlabel ndcontact -3765 -626 -3761 -616 1 gnd
rlabel metal1 -3768 -642 -3744 -637 1 gnd
rlabel polycontact -3742 -608 -3738 -604 1 clk
rlabel metal1 -3727 -588 -3693 -584 1 vdd
rlabel pdcontact -3721 -604 -3717 -594 1 vdd
rlabel ndcontact -3721 -624 -3717 -619 1 gnd
rlabel metal1 -3727 -633 -3693 -630 1 gnd
rlabel metal1 -3297 -526 -3265 -523 5 vdd
rlabel pdcontact -3291 -550 -3287 -530 1 vdd
rlabel metal1 -3297 -582 -3265 -579 1 gnd
rlabel ndcontact -3291 -574 -3287 -569 1 gnd
rlabel polycontact -3267 -563 -3263 -559 1 clk
rlabel metal1 -3245 -526 -3221 -523 5 vdd
rlabel pdcontact -3239 -550 -3235 -540 1 vdd
rlabel metal1 -3250 -603 -3216 -598 1 gnd
rlabel ndcontact -3224 -585 -3220 -575 1 gnd
rlabel polycontact -3238 -563 -3234 -559 1 clk
rlabel metal1 -3211 -526 -3187 -523 1 vdd
rlabel pdcontact -3205 -543 -3201 -533 1 vdd
rlabel ndcontact -3205 -585 -3201 -575 1 gnd
rlabel metal1 -3208 -601 -3184 -596 1 gnd
rlabel polycontact -3182 -567 -3178 -563 1 clk
rlabel metal1 -3167 -547 -3133 -543 1 vdd
rlabel pdcontact -3161 -563 -3157 -553 1 vdd
rlabel ndcontact -3161 -583 -3157 -578 1 gnd
rlabel metal1 -3167 -592 -3133 -589 1 gnd
rlabel metal1 -4276 -1626 -4244 -1623 5 vdd
rlabel pdcontact -4270 -1650 -4266 -1630 1 vdd
rlabel metal1 -4276 -1682 -4244 -1679 1 gnd
rlabel ndcontact -4270 -1674 -4266 -1669 1 gnd
rlabel polycontact -4246 -1663 -4242 -1659 1 clk
rlabel metal1 -4224 -1626 -4200 -1623 5 vdd
rlabel pdcontact -4218 -1650 -4214 -1640 1 vdd
rlabel metal1 -4229 -1703 -4195 -1698 1 gnd
rlabel ndcontact -4203 -1685 -4199 -1675 1 gnd
rlabel polycontact -4217 -1663 -4213 -1659 1 clk
rlabel metal1 -4190 -1626 -4166 -1623 1 vdd
rlabel pdcontact -4184 -1643 -4180 -1633 1 vdd
rlabel ndcontact -4184 -1685 -4180 -1675 1 gnd
rlabel metal1 -4187 -1701 -4163 -1696 1 gnd
rlabel polycontact -4161 -1667 -4157 -1663 1 clk
rlabel metal1 -4146 -1647 -4112 -1643 1 vdd
rlabel pdcontact -4140 -1663 -4136 -1653 1 vdd
rlabel ndcontact -4140 -1683 -4136 -1678 1 gnd
rlabel metal1 -4146 -1692 -4112 -1689 1 gnd
rlabel metal1 -4257 -1817 -4225 -1814 5 vdd
rlabel pdcontact -4251 -1841 -4247 -1821 1 vdd
rlabel metal1 -4257 -1873 -4225 -1870 1 gnd
rlabel ndcontact -4251 -1865 -4247 -1860 1 gnd
rlabel polycontact -4227 -1854 -4223 -1850 1 clk
rlabel metal1 -4205 -1817 -4181 -1814 5 vdd
rlabel pdcontact -4199 -1841 -4195 -1831 1 vdd
rlabel metal1 -4210 -1894 -4176 -1889 1 gnd
rlabel ndcontact -4184 -1876 -4180 -1866 1 gnd
rlabel polycontact -4198 -1854 -4194 -1850 1 clk
rlabel metal1 -4171 -1817 -4147 -1814 1 vdd
rlabel pdcontact -4165 -1834 -4161 -1824 1 vdd
rlabel ndcontact -4165 -1876 -4161 -1866 1 gnd
rlabel metal1 -4168 -1892 -4144 -1887 1 gnd
rlabel polycontact -4142 -1858 -4138 -1854 1 clk
rlabel metal1 -4127 -1838 -4093 -1834 1 vdd
rlabel pdcontact -4121 -1854 -4117 -1844 1 vdd
rlabel ndcontact -4121 -1874 -4117 -1869 1 gnd
rlabel metal1 -4127 -1883 -4093 -1880 1 gnd
rlabel metal1 -3633 -1978 -3601 -1975 5 vdd
rlabel pdcontact -3627 -2002 -3623 -1982 1 vdd
rlabel metal1 -3633 -2034 -3601 -2031 1 gnd
rlabel ndcontact -3627 -2026 -3623 -2021 1 gnd
rlabel polycontact -3603 -2015 -3599 -2011 1 clk
rlabel metal1 -3581 -1978 -3557 -1975 5 vdd
rlabel pdcontact -3575 -2002 -3571 -1992 1 vdd
rlabel metal1 -3586 -2055 -3552 -2050 1 gnd
rlabel ndcontact -3560 -2037 -3556 -2027 1 gnd
rlabel polycontact -3574 -2015 -3570 -2011 1 clk
rlabel metal1 -3547 -1978 -3523 -1975 1 vdd
rlabel pdcontact -3541 -1995 -3537 -1985 1 vdd
rlabel ndcontact -3541 -2037 -3537 -2027 1 gnd
rlabel metal1 -3544 -2053 -3520 -2048 1 gnd
rlabel polycontact -3518 -2019 -3514 -2015 1 clk
rlabel metal1 -3503 -1999 -3469 -1995 1 vdd
rlabel pdcontact -3497 -2015 -3493 -2005 1 vdd
rlabel ndcontact -3497 -2035 -3493 -2030 1 gnd
rlabel metal1 -3503 -2044 -3469 -2041 1 gnd
rlabel metal1 -3334 -1969 -3302 -1966 5 vdd
rlabel pdcontact -3328 -1993 -3324 -1973 1 vdd
rlabel metal1 -3334 -2025 -3302 -2022 1 gnd
rlabel ndcontact -3328 -2017 -3324 -2012 1 gnd
rlabel polycontact -3304 -2006 -3300 -2002 1 clk
rlabel metal1 -3282 -1969 -3258 -1966 5 vdd
rlabel pdcontact -3276 -1993 -3272 -1983 1 vdd
rlabel metal1 -3287 -2046 -3253 -2041 1 gnd
rlabel ndcontact -3261 -2028 -3257 -2018 1 gnd
rlabel polycontact -3275 -2006 -3271 -2002 1 clk
rlabel metal1 -3248 -1969 -3224 -1966 1 vdd
rlabel pdcontact -3242 -1986 -3238 -1976 1 vdd
rlabel ndcontact -3242 -2028 -3238 -2018 1 gnd
rlabel metal1 -3245 -2044 -3221 -2039 1 gnd
rlabel polycontact -3219 -2010 -3215 -2006 1 clk
rlabel metal1 -3204 -1990 -3170 -1986 1 vdd
rlabel pdcontact -3198 -2006 -3194 -1996 1 vdd
rlabel ndcontact -3198 -2026 -3194 -2021 1 gnd
rlabel metal1 -3204 -2035 -3170 -2032 1 gnd
rlabel metal1 -2958 -1820 -2926 -1817 5 vdd
rlabel pdcontact -2952 -1844 -2948 -1824 1 vdd
rlabel metal1 -2958 -1876 -2926 -1873 1 gnd
rlabel ndcontact -2952 -1868 -2948 -1863 1 gnd
rlabel polycontact -2928 -1857 -2924 -1853 1 clk
rlabel metal1 -2906 -1820 -2882 -1817 5 vdd
rlabel pdcontact -2900 -1844 -2896 -1834 1 vdd
rlabel metal1 -2911 -1897 -2877 -1892 1 gnd
rlabel ndcontact -2885 -1879 -2881 -1869 1 gnd
rlabel polycontact -2899 -1857 -2895 -1853 1 clk
rlabel metal1 -2872 -1820 -2848 -1817 1 vdd
rlabel pdcontact -2866 -1837 -2862 -1827 1 vdd
rlabel ndcontact -2866 -1879 -2862 -1869 1 gnd
rlabel metal1 -2869 -1895 -2845 -1890 1 gnd
rlabel polycontact -2843 -1861 -2839 -1857 1 clk
rlabel metal1 -2828 -1841 -2794 -1837 1 vdd
rlabel pdcontact -2822 -1857 -2818 -1847 1 vdd
rlabel ndcontact -2822 -1877 -2818 -1872 1 gnd
rlabel metal1 -2828 -1886 -2794 -1883 1 gnd
rlabel metal1 -2720 -1816 -2688 -1813 5 vdd
rlabel pdcontact -2714 -1840 -2710 -1820 1 vdd
rlabel metal1 -2720 -1872 -2688 -1869 1 gnd
rlabel ndcontact -2714 -1864 -2710 -1859 1 gnd
rlabel polycontact -2690 -1853 -2686 -1849 1 clk
rlabel metal1 -2668 -1816 -2644 -1813 5 vdd
rlabel pdcontact -2662 -1840 -2658 -1830 1 vdd
rlabel metal1 -2673 -1893 -2639 -1888 1 gnd
rlabel ndcontact -2647 -1875 -2643 -1865 1 gnd
rlabel polycontact -2661 -1853 -2657 -1849 1 clk
rlabel metal1 -2634 -1816 -2610 -1813 1 vdd
rlabel pdcontact -2628 -1833 -2624 -1823 1 vdd
rlabel ndcontact -2628 -1875 -2624 -1865 1 gnd
rlabel metal1 -2631 -1891 -2607 -1886 1 gnd
rlabel polycontact -2605 -1857 -2601 -1853 1 clk
rlabel metal1 -2590 -1837 -2556 -1833 1 vdd
rlabel pdcontact -2584 -1853 -2580 -1843 1 vdd
rlabel ndcontact -2584 -1873 -2580 -1868 1 gnd
rlabel metal1 -2590 -1882 -2556 -1879 1 gnd
rlabel metal1 -2271 -1805 -2239 -1802 5 vdd
rlabel pdcontact -2265 -1829 -2261 -1809 1 vdd
rlabel metal1 -2271 -1861 -2239 -1858 1 gnd
rlabel ndcontact -2265 -1853 -2261 -1848 1 gnd
rlabel polycontact -2241 -1842 -2237 -1838 1 clk
rlabel metal1 -2219 -1805 -2195 -1802 5 vdd
rlabel pdcontact -2213 -1829 -2209 -1819 1 vdd
rlabel metal1 -2224 -1882 -2190 -1877 1 gnd
rlabel ndcontact -2198 -1864 -2194 -1854 1 gnd
rlabel polycontact -2212 -1842 -2208 -1838 1 clk
rlabel metal1 -2185 -1805 -2161 -1802 1 vdd
rlabel pdcontact -2179 -1822 -2175 -1812 1 vdd
rlabel ndcontact -2179 -1864 -2175 -1854 1 gnd
rlabel metal1 -2182 -1880 -2158 -1875 1 gnd
rlabel polycontact -2156 -1846 -2152 -1842 1 clk
rlabel metal1 -2141 -1826 -2107 -1822 1 vdd
rlabel pdcontact -2135 -1842 -2131 -1832 1 vdd
rlabel ndcontact -2135 -1862 -2131 -1857 1 gnd
rlabel metal1 -2141 -1871 -2107 -1868 1 gnd
rlabel metal1 -1954 -1798 -1922 -1795 5 vdd
rlabel pdcontact -1948 -1822 -1944 -1802 1 vdd
rlabel metal1 -1954 -1854 -1922 -1851 1 gnd
rlabel ndcontact -1948 -1846 -1944 -1841 1 gnd
rlabel polycontact -1924 -1835 -1920 -1831 1 clk
rlabel metal1 -1902 -1798 -1878 -1795 5 vdd
rlabel pdcontact -1896 -1822 -1892 -1812 1 vdd
rlabel metal1 -1907 -1875 -1873 -1870 1 gnd
rlabel ndcontact -1881 -1857 -1877 -1847 1 gnd
rlabel polycontact -1895 -1835 -1891 -1831 1 clk
rlabel metal1 -1868 -1798 -1844 -1795 1 vdd
rlabel pdcontact -1862 -1815 -1858 -1805 1 vdd
rlabel ndcontact -1862 -1857 -1858 -1847 1 gnd
rlabel metal1 -1865 -1873 -1841 -1868 1 gnd
rlabel polycontact -1839 -1839 -1835 -1835 1 clk
rlabel metal1 -1824 -1819 -1790 -1815 1 vdd
rlabel pdcontact -1818 -1835 -1814 -1825 1 vdd
rlabel ndcontact -1818 -1855 -1814 -1850 1 gnd
rlabel metal1 -1824 -1864 -1790 -1861 1 gnd
rlabel metal1 -2298 -517 -2266 -514 5 vdd
rlabel pdcontact -2292 -541 -2288 -521 1 vdd
rlabel metal1 -2298 -573 -2266 -570 1 gnd
rlabel ndcontact -2292 -565 -2288 -560 1 gnd
rlabel polycontact -2268 -554 -2264 -550 1 clk
rlabel metal1 -2246 -517 -2222 -514 5 vdd
rlabel pdcontact -2240 -541 -2236 -531 1 vdd
rlabel metal1 -2251 -594 -2217 -589 1 gnd
rlabel ndcontact -2225 -576 -2221 -566 1 gnd
rlabel polycontact -2239 -554 -2235 -550 1 clk
rlabel metal1 -2212 -517 -2188 -514 1 vdd
rlabel pdcontact -2206 -534 -2202 -524 1 vdd
rlabel ndcontact -2206 -576 -2202 -566 1 gnd
rlabel metal1 -2209 -592 -2185 -587 1 gnd
rlabel polycontact -2183 -558 -2179 -554 1 clk
rlabel metal1 -2168 -538 -2134 -534 1 vdd
rlabel pdcontact -2162 -554 -2158 -544 1 vdd
rlabel ndcontact -2162 -574 -2158 -569 1 gnd
rlabel metal1 -2168 -583 -2134 -580 1 gnd
rlabel metal1 -1668 -496 -1636 -493 5 vdd
rlabel pdcontact -1662 -520 -1658 -500 1 vdd
rlabel metal1 -1668 -552 -1636 -549 1 gnd
rlabel ndcontact -1662 -544 -1658 -539 1 gnd
rlabel polycontact -1638 -533 -1634 -529 1 clk
rlabel metal1 -1616 -496 -1592 -493 5 vdd
rlabel pdcontact -1610 -520 -1606 -510 1 vdd
rlabel metal1 -1621 -573 -1587 -568 1 gnd
rlabel ndcontact -1595 -555 -1591 -545 1 gnd
rlabel polycontact -1609 -533 -1605 -529 1 clk
rlabel metal1 -1582 -496 -1558 -493 1 vdd
rlabel pdcontact -1576 -513 -1572 -503 1 vdd
rlabel ndcontact -1576 -555 -1572 -545 1 gnd
rlabel metal1 -1579 -571 -1555 -566 1 gnd
rlabel polycontact -1553 -537 -1549 -533 1 clk
rlabel metal1 -1538 -517 -1504 -513 1 vdd
rlabel pdcontact -1532 -533 -1528 -523 1 vdd
rlabel ndcontact -1532 -553 -1528 -548 1 gnd
rlabel metal1 -1538 -562 -1504 -559 1 gnd
rlabel metal1 -1830 -1271 -1798 -1268 5 vdd
rlabel pdcontact -1824 -1295 -1820 -1275 1 vdd
rlabel metal1 -1830 -1327 -1798 -1324 1 gnd
rlabel ndcontact -1824 -1319 -1820 -1314 1 gnd
rlabel polycontact -1800 -1308 -1796 -1304 1 clk
rlabel metal1 -1778 -1271 -1754 -1268 5 vdd
rlabel pdcontact -1772 -1295 -1768 -1285 1 vdd
rlabel metal1 -1783 -1348 -1749 -1343 1 gnd
rlabel ndcontact -1757 -1330 -1753 -1320 1 gnd
rlabel polycontact -1771 -1308 -1767 -1304 1 clk
rlabel metal1 -1744 -1271 -1720 -1268 1 vdd
rlabel pdcontact -1738 -1288 -1734 -1278 1 vdd
rlabel ndcontact -1738 -1330 -1734 -1320 1 gnd
rlabel metal1 -1741 -1346 -1717 -1341 1 gnd
rlabel polycontact -1715 -1312 -1711 -1308 1 clk
rlabel metal1 -1700 -1292 -1666 -1288 1 vdd
rlabel pdcontact -1694 -1308 -1690 -1298 1 vdd
rlabel ndcontact -1694 -1328 -1690 -1323 1 gnd
rlabel metal1 -1700 -1337 -1666 -1334 1 gnd
rlabel pdiffusion -4296 -1339 -4292 -1319 1 m23c0
rlabel pdcontact -4288 -1339 -4284 -1319 1 xc0
rlabel ndcontact -4288 -1363 -4284 -1358 1 xc0
rlabel polycontact -4260 -1361 -4255 -1356 1 xc0
rlabel pdcontact -4244 -1339 -4240 -1329 1 yc0
rlabel ndcontact -4260 -1374 -4256 -1364 1 yc0
rlabel ndiffusion -4252 -1374 -4248 -1364 1 m45c0
rlabel polycontact -4217 -1361 -4213 -1357 1 yc0
rlabel ndiffusion -4210 -1374 -4206 -1364 1 m78c0
rlabel pdcontact -4210 -1332 -4206 -1322 1 c0dn
rlabel ndcontact -4202 -1374 -4198 -1364 1 c0dn
rlabel polycontact -4172 -1364 -4168 -1360 1 c0dn
rlabel pdcontact -4156 -1352 -4152 -1342 1 c0
rlabel ndcontact -4156 -1372 -4152 -1367 1 c0
rlabel metal1 -4152 -1364 -4146 -1359 1 c0
rlabel polycontact -4303 -1351 -4299 -1347 1 c01
rlabel polycontact -4269 -1662 -4265 -1658 1 b01
rlabel pdiffusion -4262 -1650 -4258 -1630 1 m23b0
rlabel pdcontact -4254 -1650 -4250 -1630 1 xb0
rlabel ndcontact -4254 -1674 -4250 -1669 1 xb0
rlabel polycontact -4226 -1672 -4221 -1667 1 xb0
rlabel pdcontact -4210 -1650 -4206 -1640 1 yb0
rlabel ndcontact -4226 -1685 -4222 -1675 1 yb0
rlabel polycontact -4183 -1672 -4179 -1668 1 yb0
rlabel ndiffusion -4218 -1685 -4214 -1675 1 m45b0
rlabel ndiffusion -4176 -1685 -4172 -1675 1 m78b0
rlabel pdcontact -4176 -1643 -4172 -1633 1 b0dn
rlabel ndcontact -4168 -1685 -4164 -1675 1 b0dn
rlabel polycontact -4138 -1675 -4134 -1671 1 b0dn
rlabel ndcontact -4122 -1683 -4118 -1678 1 b0
rlabel pdcontact -4122 -1663 -4118 -1653 1 b0
rlabel metal1 -4116 -1675 -4112 -1670 1 b0
rlabel m3contact -3858 -1675 -3851 -1670 1 b0
rlabel polycontact -4250 -1853 -4246 -1849 1 a01
rlabel pdiffusion -4243 -1841 -4239 -1821 1 m23a0
rlabel pdcontact -4235 -1841 -4231 -1821 1 xa0
rlabel ndcontact -4235 -1865 -4231 -1860 1 xa0
rlabel polycontact -4207 -1863 -4202 -1858 1 xa0
rlabel pdcontact -4191 -1841 -4187 -1831 1 ya0
rlabel ndcontact -4207 -1876 -4203 -1866 1 ya0
rlabel ndiffusion -4199 -1876 -4195 -1866 1 m45a0
rlabel polycontact -4164 -1863 -4160 -1859 1 ya0
rlabel ndiffusion -4157 -1876 -4153 -1866 1 m78a0
rlabel pdcontact -4157 -1834 -4153 -1824 1 a0dn
rlabel ndcontact -4149 -1876 -4145 -1866 1 a0dn
rlabel polycontact -4119 -1866 -4115 -1862 1 a0dn
rlabel ndcontact -4103 -1874 -4099 -1869 1 a0
rlabel pdcontact -4103 -1854 -4099 -1844 1 a0
rlabel metal1 -4097 -1866 -4091 -1861 1 a0
rlabel m3contact -3879 -1766 -3871 -1760 1 a0
rlabel polycontact -3626 -2014 -3622 -2010 1 a11
rlabel pdiffusion -3619 -2002 -3615 -1982 1 m23a11
rlabel pdcontact -3611 -2002 -3607 -1982 1 xa11
rlabel ndcontact -3611 -2026 -3607 -2021 1 xa11
rlabel polycontact -3583 -2024 -3578 -2019 1 xa11
rlabel pdcontact -3567 -2002 -3563 -1992 1 ya11
rlabel ndcontact -3583 -2037 -3579 -2027 1 ya11
rlabel ndiffusion -3575 -2037 -3571 -2027 1 m45a11
rlabel polycontact -3540 -2024 -3536 -2020 1 ya11
rlabel ndiffusion -3533 -2037 -3529 -2027 1 m78a11
rlabel ndcontact -3525 -2037 -3521 -2027 1 a1dn
rlabel pdcontact -3533 -1995 -3529 -1985 1 a1dn
rlabel polycontact -3495 -2027 -3491 -2023 1 a1dn
rlabel metal1 -3475 -2027 -3469 -2022 1 a1
rlabel m3contact -3516 -1779 -3509 -1774 1 a1
rlabel pdiffusion -3320 -1993 -3316 -1973 1 m23b1
rlabel pdcontact -3312 -1993 -3308 -1973 1 xb1
rlabel ndcontact -3312 -2017 -3308 -2012 1 xb1
rlabel polycontact -3284 -2015 -3279 -2010 1 xb1
rlabel ndcontact -3284 -2028 -3280 -2018 1 yb1
rlabel pdcontact -3268 -1993 -3264 -1983 1 yb1
rlabel polycontact -3241 -2015 -3237 -2011 1 yb1
rlabel ndiffusion -3276 -2028 -3272 -2018 1 m45b1
rlabel ndiffusion -3234 -2028 -3230 -2018 1 m78b1
rlabel pdcontact -3234 -1986 -3230 -1976 1 b1dn
rlabel ndcontact -3226 -2028 -3222 -2018 1 b1dn
rlabel polycontact -3196 -2018 -3192 -2014 1 b1dn
rlabel pdcontact -3479 -2015 -3475 -2005 1 a1
rlabel ndcontact -3479 -2035 -3475 -2030 1 a1
rlabel ndcontact -3180 -2026 -3176 -2021 1 b1
rlabel pdcontact -3180 -2006 -3176 -1996 1 b1
rlabel metal1 -3174 -2018 -3169 -2013 1 b1
rlabel polycontact -2951 -1856 -2947 -1852 1 a21
rlabel pdiffusion -2944 -1844 -2940 -1824 1 m23a2
rlabel pdcontact -2936 -1844 -2932 -1824 1 xa2
rlabel ndcontact -2936 -1868 -2932 -1863 1 xa2
rlabel polycontact -2908 -1866 -2903 -1861 1 xa2
rlabel pdcontact -2892 -1844 -2888 -1834 1 ya2
rlabel ndcontact -2908 -1879 -2904 -1869 1 ya2
rlabel ndiffusion -2900 -1879 -2896 -1869 1 m45a2
rlabel polycontact -2865 -1866 -2861 -1862 1 ya2
rlabel ndiffusion -2858 -1879 -2854 -1869 1 m78a2
rlabel ndcontact -2850 -1879 -2846 -1869 1 a2dn
rlabel pdcontact -2858 -1837 -2854 -1827 1 a2dn
rlabel polycontact -2820 -1869 -2816 -1865 1 a2dn
rlabel pdcontact -2804 -1857 -2800 -1847 1 a2
rlabel ndcontact -2804 -1877 -2800 -1872 1 a2
rlabel metal1 -2798 -1869 -2794 -1864 1 a2
rlabel m3contact -2972 -1686 -2967 -1680 1 a2
rlabel pdiffusion -2706 -1840 -2702 -1820 1 m23b2
rlabel pdcontact -2698 -1840 -2694 -1820 1 xb2
rlabel ndcontact -2698 -1864 -2694 -1859 1 xb2
rlabel polycontact -2670 -1862 -2665 -1857 1 xb2
rlabel ndcontact -2670 -1875 -2666 -1865 1 yb2
rlabel ndiffusion -2662 -1875 -2658 -1865 1 m45b2
rlabel pdcontact -2654 -1840 -2650 -1830 1 yb2
rlabel polycontact -2627 -1862 -2623 -1858 1 yb2
rlabel ndiffusion -2620 -1875 -2616 -1865 1 m78b2
rlabel ndcontact -2612 -1875 -2608 -1865 1 b2dn
rlabel pdcontact -2620 -1833 -2616 -1823 1 b2dn
rlabel polycontact -2582 -1865 -2578 -1861 1 b2dn
rlabel pdcontact -2566 -1853 -2562 -1843 1 b2
rlabel ndcontact -2566 -1873 -2562 -1868 1 b2
rlabel metal1 -2560 -1865 -2556 -1860 1 b2
rlabel metal2 -2837 -1740 -2832 -1734 1 b2
rlabel polycontact -2264 -1841 -2260 -1837 1 a31
rlabel pdiffusion -2257 -1829 -2253 -1809 1 m23a3
rlabel pdcontact -2249 -1829 -2245 -1809 1 xa3
rlabel ndcontact -2249 -1853 -2245 -1848 1 xa3
rlabel polycontact -2221 -1851 -2216 -1846 1 xa3
rlabel ndcontact -2221 -1864 -2217 -1854 1 ya3
rlabel ndiffusion -2213 -1864 -2209 -1854 1 m45a3
rlabel pdcontact -2205 -1829 -2201 -1819 1 ya3
rlabel ndiffusion -2171 -1864 -2167 -1854 1 m78a3
rlabel ndcontact -2163 -1864 -2159 -1854 1 a3dn
rlabel pdcontact -2171 -1822 -2167 -1812 1 a3dn
rlabel polycontact -2178 -1851 -2174 -1847 1 ya3
rlabel polycontact -2133 -1854 -2129 -1850 1 a3dn
rlabel ndcontact -2117 -1862 -2113 -1857 1 a3
rlabel pdcontact -2117 -1842 -2113 -1832 1 a3
rlabel m3contact -2253 -1591 -2248 -1583 1 a3
rlabel polycontact -2181 -1747 -2177 -1743 1 b3
rlabel pdiffusion -1940 -1822 -1936 -1802 1 m23b3
rlabel pdcontact -1932 -1822 -1928 -1802 1 xb3
rlabel ndcontact -1932 -1846 -1928 -1841 1 xb3
rlabel polycontact -1904 -1844 -1899 -1839 1 xb3
rlabel ndcontact -1904 -1857 -1900 -1847 1 yb3
rlabel pdcontact -1888 -1822 -1884 -1812 1 yb3
rlabel polycontact -1861 -1844 -1857 -1840 1 yb3
rlabel ndiffusion -1896 -1857 -1892 -1847 1 m45b3
rlabel ndiffusion -1854 -1857 -1850 -1847 1 m78b3
rlabel ndcontact -1846 -1857 -1842 -1847 1 b3dn
rlabel pdcontact -1854 -1815 -1850 -1805 1 b3dn
rlabel polycontact -1816 -1847 -1812 -1843 1 b3dn
rlabel ndcontact -1800 -1855 -1796 -1850 1 b3
rlabel pdcontact -1800 -1835 -1796 -1825 1 b3
rlabel m3contact -2167 -1716 -2162 -1711 1 b3
rlabel polycontact -3850 -603 -3846 -599 1 s0
rlabel ndcontact -3835 -615 -3831 -610 1 xs0
rlabel pdiffusion -3843 -591 -3839 -571 1 m23s0
rlabel pdcontact -3835 -591 -3831 -571 1 xs0
rlabel polycontact -3807 -613 -3802 -608 1 xs0
rlabel ndcontact -3807 -626 -3803 -616 1 ys0
rlabel pdcontact -3791 -591 -3787 -581 1 ys0
rlabel ndiffusion -3799 -626 -3795 -616 1 m45s0
rlabel polycontact -3764 -613 -3760 -609 1 ys0
rlabel ndcontact -3749 -626 -3745 -616 1 s0dn
rlabel pdcontact -3757 -584 -3753 -574 1 s0dn
rlabel polycontact -3719 -616 -3715 -612 1 s0dn
rlabel metal1 -3697 -616 -3690 -611 1 s0f
rlabel ndcontact -3703 -624 -3699 -619 1 s0f
rlabel pdcontact -3703 -604 -3699 -594 1 s0f
rlabel pdiffusion -3283 -550 -3279 -530 1 m23s1
rlabel pdcontact -3275 -550 -3271 -530 1 xs1
rlabel ndcontact -3275 -574 -3271 -569 1 xs1
rlabel polycontact -3247 -572 -3242 -567 1 xs1
rlabel polycontact -3290 -562 -3286 -558 1 s1
rlabel ndcontact -3247 -585 -3243 -575 1 ys1
rlabel ndiffusion -3239 -585 -3235 -575 1 m45s1
rlabel pdcontact -3231 -550 -3227 -540 1 ys1
rlabel polycontact -3204 -572 -3200 -568 1 ys1
rlabel ndiffusion -3197 -585 -3193 -575 1 m78s1
rlabel ndcontact -3189 -585 -3185 -575 1 s1dn
rlabel pdcontact -3197 -543 -3193 -533 1 s1dn
rlabel polycontact -3159 -575 -3155 -571 1 s1dn
rlabel pdcontact -3143 -563 -3139 -553 1 s1f
rlabel ndcontact -3143 -583 -3139 -578 1 s1f
rlabel metal1 -3137 -575 -3133 -571 1 s1f
rlabel polycontact -2291 -553 -2287 -549 1 s2
rlabel ndcontact -2276 -565 -2272 -560 1 xs2
rlabel pdcontact -2276 -541 -2272 -521 1 xs2
rlabel pdiffusion -2284 -541 -2280 -521 1 m23s2
rlabel polycontact -2248 -563 -2243 -558 1 xs2
rlabel ndcontact -2248 -576 -2244 -566 1 ys2
rlabel ndiffusion -2240 -576 -2236 -566 1 m45s2
rlabel polycontact -2205 -563 -2201 -559 1 ys2
rlabel ndiffusion -2198 -576 -2194 -566 1 m78s2
rlabel ndcontact -2190 -576 -2186 -566 1 s2dn
rlabel pdcontact -2198 -534 -2194 -524 1 s2dn
rlabel polycontact -2160 -566 -2156 -562 1 s2dn
rlabel ndcontact -2144 -574 -2140 -569 1 s2f
rlabel pdcontact -2144 -554 -2140 -544 1 s2f
rlabel metal1 -2138 -566 -2134 -562 1 s2f
rlabel polycontact -1661 -532 -1657 -528 1 s3
rlabel ndcontact -1646 -544 -1642 -539 1 xs3
rlabel pdcontact -1646 -520 -1642 -500 1 xs3
rlabel polycontact -1618 -542 -1613 -537 1 xs3
rlabel ndcontact -1618 -555 -1614 -545 1 ys3
rlabel pdcontact -1602 -520 -1598 -510 1 ys3
rlabel ndiffusion -1610 -555 -1606 -545 1 m45s3
rlabel polycontact -1575 -542 -1571 -538 1 ys3
rlabel ndiffusion -1568 -555 -1564 -545 1 m78s3
rlabel ndcontact -1560 -555 -1556 -545 1 s3dn
rlabel pdcontact -1568 -513 -1564 -503 1 s3dn
rlabel polycontact -1530 -545 -1526 -541 1 s3dn
rlabel ndcontact -1514 -553 -1510 -548 1 s3f
rlabel pdcontact -1514 -533 -1510 -523 1 s3f
rlabel metal1 -1508 -545 -1504 -541 7 s3f
rlabel metal1 -1670 -1320 -1666 -1316 1 c4f
rlabel ndcontact -1676 -1328 -1672 -1323 1 c4f
rlabel pdcontact -1676 -1308 -1672 -1298 1 c4f
rlabel polycontact -1692 -1320 -1688 -1316 1 c4dn
rlabel ndcontact -1722 -1330 -1718 -1320 1 c4dn
rlabel pdcontact -1730 -1288 -1726 -1278 1 c4dn
rlabel ndiffusion -1730 -1330 -1726 -1320 1 m78c4
rlabel ndiffusion -1772 -1330 -1768 -1320 1 m45c4
rlabel ndcontact -1780 -1330 -1776 -1320 1 yc4
rlabel pdcontact -1764 -1295 -1760 -1285 1 yc4
rlabel polycontact -1737 -1317 -1733 -1313 1 yc4
rlabel polycontact -1780 -1317 -1775 -1312 1 xc4
rlabel ndcontact -1808 -1319 -1804 -1314 1 xc4
rlabel pdcontact -1808 -1295 -1804 -1275 1 xc4
rlabel pdiffusion -1816 -1295 -1812 -1275 1 m23c4
rlabel polycontact -1823 -1307 -1819 -1303 1 c4
rlabel ndiffusion -3757 -626 -3753 -616 1 m78s0
rlabel pdiffusion -1654 -520 -1650 -500 1 m23s3
rlabel pdcontact -2232 -541 -2228 -531 1 ys2
rlabel metal1 -2111 -1854 -2106 -1849 1 a3
rlabel metal1 -1794 -1847 -1781 -1842 1 b3
rlabel metal1 -3642 -1532 -3629 -1527 1 c1
rlabel polycontact -3327 -2005 -3323 -2001 1 b11
rlabel polycontact -2713 -1852 -2709 -1848 1 b21
rlabel polycontact -1947 -1834 -1943 -1830 1 b31
<< end >>
