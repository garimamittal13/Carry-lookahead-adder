magic
tech scmos
timestamp 1732060801
<< nwell >>
rect 1123 3824 1157 3850
rect 1169 3834 1203 3859
rect 1217 3831 1251 3857
rect 1844 3850 1878 3876
rect 1890 3860 1924 3885
rect 1938 3857 1972 3883
rect 2466 3868 2500 3894
rect 2512 3878 2546 3903
rect 2560 3875 2594 3901
rect 1123 3768 1157 3794
rect 1171 3768 1205 3793
rect 1219 3765 1253 3791
rect 1277 3788 1311 3826
rect 1326 3791 1360 3817
rect 1844 3794 1878 3820
rect 1892 3794 1926 3819
rect 1940 3791 1974 3817
rect 1998 3814 2032 3852
rect 2047 3817 2081 3843
rect 2466 3812 2500 3838
rect 2514 3812 2548 3837
rect 2562 3809 2596 3835
rect 2620 3832 2654 3870
rect 2669 3835 2703 3861
rect 578 3578 612 3604
rect 624 3588 658 3613
rect 672 3585 706 3611
rect 578 3522 612 3548
rect 626 3522 660 3547
rect 674 3519 708 3545
rect 732 3542 766 3580
rect 781 3545 815 3571
rect 1964 3482 1998 3507
rect 2012 3479 2046 3505
rect 2103 3423 2137 3461
rect 2152 3426 2186 3452
rect 1963 3359 1997 3384
rect 2011 3356 2045 3382
rect 1479 3326 1513 3351
rect 1527 3323 1561 3349
rect 1611 3278 1645 3316
rect 1660 3281 1694 3307
rect 2279 3303 2313 3341
rect 2328 3306 2362 3332
rect 2464 3312 2498 3350
rect 2513 3315 2547 3341
rect 907 3209 941 3234
rect 955 3206 989 3232
rect 1478 3220 1512 3245
rect 1526 3217 1560 3243
rect 1727 3239 1761 3277
rect 1776 3242 1810 3268
rect 1968 3236 2002 3261
rect 2016 3233 2050 3259
rect 1033 3135 1067 3173
rect 1082 3138 1116 3164
rect 1148 3145 1182 3183
rect 1615 3176 1649 3214
rect 1664 3179 1698 3205
rect 2102 3179 2136 3217
rect 2151 3182 2185 3208
rect 1197 3148 1231 3174
rect 573 3091 607 3116
rect 621 3088 655 3114
rect 677 3087 711 3125
rect 726 3090 760 3116
rect 912 3100 946 3125
rect 1482 3123 1516 3148
rect 960 3097 994 3123
rect 1530 3120 1564 3146
rect 1967 3108 2001 3133
rect 2015 3105 2049 3131
rect 576 2988 610 3014
rect 622 2998 656 3023
rect 670 2995 704 3021
rect 928 2990 962 3016
rect 974 3000 1008 3025
rect 1022 2997 1056 3023
rect 576 2932 610 2958
rect 624 2932 658 2957
rect 672 2929 706 2955
rect 730 2952 764 2990
rect 779 2955 813 2981
rect 928 2934 962 2960
rect 976 2934 1010 2959
rect 1024 2931 1058 2957
rect 1082 2954 1116 2992
rect 1489 2990 1523 3016
rect 1535 3000 1569 3025
rect 1583 2997 1617 3023
rect 2164 3009 2198 3035
rect 2210 3019 2244 3044
rect 2258 3016 2292 3042
rect 1131 2957 1165 2983
rect 1489 2934 1523 2960
rect 1537 2934 1571 2959
rect 1585 2931 1619 2957
rect 1643 2954 1677 2992
rect 1692 2957 1726 2983
rect 2164 2953 2198 2979
rect 2212 2953 2246 2978
rect 2260 2950 2294 2976
rect 2318 2973 2352 3011
rect 2367 2976 2401 3002
rect 2199 2874 2233 2899
rect 2247 2871 2281 2897
rect 592 2823 626 2848
rect 640 2820 674 2846
rect 979 2843 1013 2868
rect 1027 2840 1061 2866
rect 1529 2844 1563 2869
rect 1577 2841 1611 2867
<< ntransistor >>
rect 2478 3854 2480 3859
rect 2523 3855 2525 3865
rect 2533 3855 2535 3865
rect 2572 3861 2574 3866
rect 1856 3836 1858 3841
rect 1901 3837 1903 3847
rect 1911 3837 1913 3847
rect 1950 3843 1952 3848
rect 1135 3810 1137 3815
rect 1180 3811 1182 3821
rect 1190 3811 1192 3821
rect 1229 3817 1231 3822
rect 1135 3754 1137 3759
rect 1338 3777 1340 3782
rect 1856 3780 1858 3785
rect 2059 3803 2061 3808
rect 2009 3795 2011 3800
rect 2019 3795 2021 3800
rect 2478 3798 2480 3803
rect 2681 3821 2683 3826
rect 2631 3813 2633 3818
rect 2641 3813 2643 3818
rect 2525 3789 2527 3799
rect 2535 3789 2537 3799
rect 2574 3795 2576 3800
rect 1288 3769 1290 3774
rect 1298 3769 1300 3774
rect 1903 3771 1905 3781
rect 1913 3771 1915 3781
rect 1952 3777 1954 3782
rect 1182 3745 1184 3755
rect 1192 3745 1194 3755
rect 1231 3751 1233 3756
rect 590 3564 592 3569
rect 635 3565 637 3575
rect 645 3565 647 3575
rect 684 3571 686 3576
rect 590 3508 592 3513
rect 793 3531 795 3536
rect 743 3523 745 3528
rect 753 3523 755 3528
rect 637 3499 639 3509
rect 647 3499 649 3509
rect 686 3505 688 3510
rect 1975 3459 1977 3469
rect 1985 3459 1987 3469
rect 2024 3465 2026 3470
rect 2164 3412 2166 3417
rect 2114 3404 2116 3409
rect 2124 3404 2126 3409
rect 1974 3336 1976 3346
rect 1984 3336 1986 3346
rect 2023 3342 2025 3347
rect 1490 3303 1492 3313
rect 1500 3303 1502 3313
rect 1539 3309 1541 3314
rect 2525 3301 2527 3306
rect 2340 3292 2342 3297
rect 2475 3293 2477 3298
rect 2485 3293 2487 3298
rect 2290 3284 2292 3289
rect 2300 3284 2302 3289
rect 1672 3267 1674 3272
rect 1622 3259 1624 3264
rect 1632 3259 1634 3264
rect 1788 3228 1790 3233
rect 1738 3220 1740 3225
rect 1748 3220 1750 3225
rect 1979 3213 1981 3223
rect 1989 3213 1991 3223
rect 2028 3219 2030 3224
rect 1489 3197 1491 3207
rect 1499 3197 1501 3207
rect 1538 3203 1540 3208
rect 918 3186 920 3196
rect 928 3186 930 3196
rect 967 3192 969 3197
rect 1676 3165 1678 3170
rect 2163 3168 2165 3173
rect 1626 3157 1628 3162
rect 1636 3157 1638 3162
rect 2113 3160 2115 3165
rect 2123 3160 2125 3165
rect 1209 3134 1211 3139
rect 1094 3124 1096 3129
rect 1159 3126 1161 3131
rect 1169 3126 1171 3131
rect 1044 3116 1046 3121
rect 1054 3116 1056 3121
rect 584 3068 586 3078
rect 594 3068 596 3078
rect 633 3074 635 3079
rect 1493 3100 1495 3110
rect 1503 3100 1505 3110
rect 1542 3106 1544 3111
rect 738 3076 740 3081
rect 923 3077 925 3087
rect 933 3077 935 3087
rect 972 3083 974 3088
rect 1978 3085 1980 3095
rect 1988 3085 1990 3095
rect 2027 3091 2029 3096
rect 688 3068 690 3073
rect 698 3068 700 3073
rect 588 2974 590 2979
rect 633 2975 635 2985
rect 643 2975 645 2985
rect 682 2981 684 2986
rect 940 2976 942 2981
rect 985 2977 987 2987
rect 995 2977 997 2987
rect 1034 2983 1036 2988
rect 2176 2995 2178 3000
rect 2221 2996 2223 3006
rect 2231 2996 2233 3006
rect 2270 3002 2272 3007
rect 588 2918 590 2923
rect 1501 2976 1503 2981
rect 1546 2977 1548 2987
rect 1556 2977 1558 2987
rect 1595 2983 1597 2988
rect 791 2941 793 2946
rect 741 2933 743 2938
rect 751 2933 753 2938
rect 940 2920 942 2925
rect 1143 2943 1145 2948
rect 1093 2935 1095 2940
rect 1103 2935 1105 2940
rect 635 2909 637 2919
rect 645 2909 647 2919
rect 684 2915 686 2920
rect 987 2911 989 2921
rect 997 2911 999 2921
rect 1036 2917 1038 2922
rect 1501 2920 1503 2925
rect 1704 2943 1706 2948
rect 1654 2935 1656 2940
rect 1664 2935 1666 2940
rect 2176 2939 2178 2944
rect 2379 2962 2381 2967
rect 2329 2954 2331 2959
rect 2339 2954 2341 2959
rect 2223 2930 2225 2940
rect 2233 2930 2235 2940
rect 2272 2936 2274 2941
rect 1548 2911 1550 2921
rect 1558 2911 1560 2921
rect 1597 2917 1599 2922
rect 2210 2851 2212 2861
rect 2220 2851 2222 2861
rect 2259 2857 2261 2862
rect 990 2820 992 2830
rect 1000 2820 1002 2830
rect 1039 2826 1041 2831
rect 1540 2821 1542 2831
rect 1550 2821 1552 2831
rect 1589 2827 1591 2832
rect 603 2800 605 2810
rect 613 2800 615 2810
rect 652 2806 654 2811
<< ptransistor >>
rect 2523 3884 2525 3894
rect 2533 3884 2535 3894
rect 1901 3866 1903 3876
rect 1911 3866 1913 3876
rect 2478 3874 2480 3884
rect 1856 3856 1858 3866
rect 1180 3840 1182 3850
rect 1190 3840 1192 3850
rect 1135 3830 1137 3840
rect 1229 3837 1231 3847
rect 1950 3863 1952 3873
rect 2572 3881 2574 3891
rect 2009 3820 2011 3840
rect 2019 3820 2021 3840
rect 2631 3838 2633 3858
rect 2641 3838 2643 3858
rect 2681 3841 2683 3851
rect 2059 3823 2061 3833
rect 1288 3794 1290 3814
rect 1298 3794 1300 3814
rect 1338 3797 1340 3807
rect 1856 3800 1858 3810
rect 1903 3800 1905 3810
rect 1913 3800 1915 3810
rect 1135 3774 1137 3784
rect 1182 3774 1184 3784
rect 1192 3774 1194 3784
rect 1231 3771 1233 3781
rect 1952 3797 1954 3807
rect 2478 3818 2480 3828
rect 2525 3818 2527 3828
rect 2535 3818 2537 3828
rect 2574 3815 2576 3825
rect 635 3594 637 3604
rect 645 3594 647 3604
rect 590 3584 592 3594
rect 684 3591 686 3601
rect 743 3548 745 3568
rect 753 3548 755 3568
rect 793 3551 795 3561
rect 590 3528 592 3538
rect 637 3528 639 3538
rect 647 3528 649 3538
rect 686 3525 688 3535
rect 1975 3488 1977 3498
rect 1985 3488 1987 3498
rect 2024 3485 2026 3495
rect 2114 3429 2116 3449
rect 2124 3429 2126 3449
rect 2164 3432 2166 3442
rect 1974 3365 1976 3375
rect 1984 3365 1986 3375
rect 2023 3362 2025 3372
rect 1490 3332 1492 3342
rect 1500 3332 1502 3342
rect 1539 3329 1541 3339
rect 2290 3309 2292 3329
rect 2300 3309 2302 3329
rect 2340 3312 2342 3322
rect 2475 3318 2477 3338
rect 2485 3318 2487 3338
rect 2525 3321 2527 3331
rect 1622 3284 1624 3304
rect 1632 3284 1634 3304
rect 1672 3287 1674 3297
rect 1738 3245 1740 3265
rect 1748 3245 1750 3265
rect 1788 3248 1790 3258
rect 1489 3226 1491 3236
rect 1499 3226 1501 3236
rect 918 3215 920 3225
rect 928 3215 930 3225
rect 967 3212 969 3222
rect 1538 3223 1540 3233
rect 1979 3242 1981 3252
rect 1989 3242 1991 3252
rect 2028 3239 2030 3249
rect 1626 3182 1628 3202
rect 1636 3182 1638 3202
rect 1676 3185 1678 3195
rect 2113 3185 2115 3205
rect 2123 3185 2125 3205
rect 2163 3188 2165 3198
rect 1044 3141 1046 3161
rect 1054 3141 1056 3161
rect 1094 3144 1096 3154
rect 1159 3151 1161 3171
rect 1169 3151 1171 3171
rect 1209 3154 1211 3164
rect 1493 3129 1495 3139
rect 1503 3129 1505 3139
rect 584 3097 586 3107
rect 594 3097 596 3107
rect 633 3094 635 3104
rect 688 3093 690 3113
rect 698 3093 700 3113
rect 923 3106 925 3116
rect 933 3106 935 3116
rect 738 3096 740 3106
rect 972 3103 974 3113
rect 1542 3126 1544 3136
rect 1978 3114 1980 3124
rect 1988 3114 1990 3124
rect 2027 3111 2029 3121
rect 2221 3025 2223 3035
rect 2231 3025 2233 3035
rect 633 3004 635 3014
rect 643 3004 645 3014
rect 588 2994 590 3004
rect 682 3001 684 3011
rect 985 3006 987 3016
rect 995 3006 997 3016
rect 940 2996 942 3006
rect 1034 3003 1036 3013
rect 1546 3006 1548 3016
rect 1556 3006 1558 3016
rect 2176 3015 2178 3025
rect 1501 2996 1503 3006
rect 741 2958 743 2978
rect 751 2958 753 2978
rect 1595 3003 1597 3013
rect 2270 3022 2272 3032
rect 791 2961 793 2971
rect 588 2938 590 2948
rect 635 2938 637 2948
rect 645 2938 647 2948
rect 684 2935 686 2945
rect 1093 2960 1095 2980
rect 1103 2960 1105 2980
rect 1143 2963 1145 2973
rect 940 2940 942 2950
rect 987 2940 989 2950
rect 997 2940 999 2950
rect 1036 2937 1038 2947
rect 1654 2960 1656 2980
rect 1664 2960 1666 2980
rect 2329 2979 2331 2999
rect 2339 2979 2341 2999
rect 2379 2982 2381 2992
rect 1704 2963 1706 2973
rect 1501 2940 1503 2950
rect 1548 2940 1550 2950
rect 1558 2940 1560 2950
rect 1597 2937 1599 2947
rect 2176 2959 2178 2969
rect 2223 2959 2225 2969
rect 2233 2959 2235 2969
rect 2272 2956 2274 2966
rect 2210 2880 2212 2890
rect 2220 2880 2222 2890
rect 2259 2877 2261 2887
rect 990 2849 992 2859
rect 1000 2849 1002 2859
rect 603 2829 605 2839
rect 613 2829 615 2839
rect 652 2826 654 2836
rect 1039 2846 1041 2856
rect 1540 2850 1542 2860
rect 1550 2850 1552 2860
rect 1589 2847 1591 2857
<< ndiffusion >>
rect 2476 3854 2478 3859
rect 2480 3854 2490 3859
rect 2522 3855 2523 3865
rect 2525 3855 2533 3865
rect 2535 3855 2536 3865
rect 2570 3861 2572 3866
rect 2574 3861 2584 3866
rect 1854 3836 1856 3841
rect 1858 3836 1868 3841
rect 1900 3837 1901 3847
rect 1903 3837 1911 3847
rect 1913 3837 1914 3847
rect 1948 3843 1950 3848
rect 1952 3843 1962 3848
rect 1133 3810 1135 3815
rect 1137 3810 1147 3815
rect 1179 3811 1180 3821
rect 1182 3811 1190 3821
rect 1192 3811 1193 3821
rect 1227 3817 1229 3822
rect 1231 3817 1241 3822
rect 1133 3754 1135 3759
rect 1137 3754 1147 3759
rect 1336 3777 1338 3782
rect 1340 3777 1350 3782
rect 1854 3780 1856 3785
rect 1858 3780 1868 3785
rect 2057 3803 2059 3808
rect 2061 3803 2071 3808
rect 2008 3795 2009 3800
rect 2011 3795 2012 3800
rect 2018 3795 2019 3800
rect 2021 3795 2022 3800
rect 2476 3798 2478 3803
rect 2480 3798 2490 3803
rect 2679 3821 2681 3826
rect 2683 3821 2693 3826
rect 2630 3813 2631 3818
rect 2633 3813 2634 3818
rect 2640 3813 2641 3818
rect 2643 3813 2644 3818
rect 2524 3789 2525 3799
rect 2527 3789 2535 3799
rect 2537 3789 2538 3799
rect 2572 3795 2574 3800
rect 2576 3795 2586 3800
rect 1287 3769 1288 3774
rect 1290 3769 1291 3774
rect 1297 3769 1298 3774
rect 1300 3769 1301 3774
rect 1902 3771 1903 3781
rect 1905 3771 1913 3781
rect 1915 3771 1916 3781
rect 1950 3777 1952 3782
rect 1954 3777 1964 3782
rect 1181 3745 1182 3755
rect 1184 3745 1192 3755
rect 1194 3745 1195 3755
rect 1229 3751 1231 3756
rect 1233 3751 1243 3756
rect 588 3564 590 3569
rect 592 3564 602 3569
rect 634 3565 635 3575
rect 637 3565 645 3575
rect 647 3565 648 3575
rect 682 3571 684 3576
rect 686 3571 696 3576
rect 588 3508 590 3513
rect 592 3508 602 3513
rect 791 3531 793 3536
rect 795 3531 805 3536
rect 742 3523 743 3528
rect 745 3523 746 3528
rect 752 3523 753 3528
rect 755 3523 756 3528
rect 636 3499 637 3509
rect 639 3499 647 3509
rect 649 3499 650 3509
rect 684 3505 686 3510
rect 688 3505 698 3510
rect 1974 3459 1975 3469
rect 1977 3459 1985 3469
rect 1987 3459 1988 3469
rect 2022 3465 2024 3470
rect 2026 3465 2036 3470
rect 2162 3412 2164 3417
rect 2166 3412 2176 3417
rect 2113 3404 2114 3409
rect 2116 3404 2117 3409
rect 2123 3404 2124 3409
rect 2126 3404 2127 3409
rect 1973 3336 1974 3346
rect 1976 3336 1984 3346
rect 1986 3336 1987 3346
rect 2021 3342 2023 3347
rect 2025 3342 2035 3347
rect 1489 3303 1490 3313
rect 1492 3303 1500 3313
rect 1502 3303 1503 3313
rect 1537 3309 1539 3314
rect 1541 3309 1551 3314
rect 2523 3301 2525 3306
rect 2527 3301 2537 3306
rect 2338 3292 2340 3297
rect 2342 3292 2352 3297
rect 2474 3293 2475 3298
rect 2477 3293 2478 3298
rect 2484 3293 2485 3298
rect 2487 3293 2488 3298
rect 2289 3284 2290 3289
rect 2292 3284 2293 3289
rect 2299 3284 2300 3289
rect 2302 3284 2303 3289
rect 1670 3267 1672 3272
rect 1674 3267 1684 3272
rect 1621 3259 1622 3264
rect 1624 3259 1625 3264
rect 1631 3259 1632 3264
rect 1634 3259 1635 3264
rect 1786 3228 1788 3233
rect 1790 3228 1800 3233
rect 1737 3220 1738 3225
rect 1740 3220 1741 3225
rect 1747 3220 1748 3225
rect 1750 3220 1751 3225
rect 1978 3213 1979 3223
rect 1981 3213 1989 3223
rect 1991 3213 1992 3223
rect 2026 3219 2028 3224
rect 2030 3219 2040 3224
rect 1488 3197 1489 3207
rect 1491 3197 1499 3207
rect 1501 3197 1502 3207
rect 1536 3203 1538 3208
rect 1540 3203 1550 3208
rect 917 3186 918 3196
rect 920 3186 928 3196
rect 930 3186 931 3196
rect 965 3192 967 3197
rect 969 3192 979 3197
rect 1674 3165 1676 3170
rect 1678 3165 1688 3170
rect 2161 3168 2163 3173
rect 2165 3168 2175 3173
rect 1625 3157 1626 3162
rect 1628 3157 1629 3162
rect 1635 3157 1636 3162
rect 1638 3157 1639 3162
rect 2112 3160 2113 3165
rect 2115 3160 2116 3165
rect 2122 3160 2123 3165
rect 2125 3160 2126 3165
rect 1207 3134 1209 3139
rect 1211 3134 1221 3139
rect 1092 3124 1094 3129
rect 1096 3124 1106 3129
rect 1158 3126 1159 3131
rect 1161 3126 1162 3131
rect 1168 3126 1169 3131
rect 1171 3126 1172 3131
rect 1043 3116 1044 3121
rect 1046 3116 1047 3121
rect 1053 3116 1054 3121
rect 1056 3116 1057 3121
rect 583 3068 584 3078
rect 586 3068 594 3078
rect 596 3068 597 3078
rect 631 3074 633 3079
rect 635 3074 645 3079
rect 1492 3100 1493 3110
rect 1495 3100 1503 3110
rect 1505 3100 1506 3110
rect 1540 3106 1542 3111
rect 1544 3106 1554 3111
rect 736 3076 738 3081
rect 740 3076 750 3081
rect 922 3077 923 3087
rect 925 3077 933 3087
rect 935 3077 936 3087
rect 970 3083 972 3088
rect 974 3083 984 3088
rect 1977 3085 1978 3095
rect 1980 3085 1988 3095
rect 1990 3085 1991 3095
rect 2025 3091 2027 3096
rect 2029 3091 2039 3096
rect 687 3068 688 3073
rect 690 3068 691 3073
rect 697 3068 698 3073
rect 700 3068 701 3073
rect 586 2974 588 2979
rect 590 2974 600 2979
rect 632 2975 633 2985
rect 635 2975 643 2985
rect 645 2975 646 2985
rect 680 2981 682 2986
rect 684 2981 694 2986
rect 938 2976 940 2981
rect 942 2976 952 2981
rect 984 2977 985 2987
rect 987 2977 995 2987
rect 997 2977 998 2987
rect 1032 2983 1034 2988
rect 1036 2983 1046 2988
rect 2174 2995 2176 3000
rect 2178 2995 2188 3000
rect 2220 2996 2221 3006
rect 2223 2996 2231 3006
rect 2233 2996 2234 3006
rect 2268 3002 2270 3007
rect 2272 3002 2282 3007
rect 586 2918 588 2923
rect 590 2918 600 2923
rect 1499 2976 1501 2981
rect 1503 2976 1513 2981
rect 1545 2977 1546 2987
rect 1548 2977 1556 2987
rect 1558 2977 1559 2987
rect 1593 2983 1595 2988
rect 1597 2983 1607 2988
rect 789 2941 791 2946
rect 793 2941 803 2946
rect 740 2933 741 2938
rect 743 2933 744 2938
rect 750 2933 751 2938
rect 753 2933 754 2938
rect 938 2920 940 2925
rect 942 2920 952 2925
rect 1141 2943 1143 2948
rect 1145 2943 1155 2948
rect 1092 2935 1093 2940
rect 1095 2935 1096 2940
rect 1102 2935 1103 2940
rect 1105 2935 1106 2940
rect 634 2909 635 2919
rect 637 2909 645 2919
rect 647 2909 648 2919
rect 682 2915 684 2920
rect 686 2915 696 2920
rect 986 2911 987 2921
rect 989 2911 997 2921
rect 999 2911 1000 2921
rect 1034 2917 1036 2922
rect 1038 2917 1048 2922
rect 1499 2920 1501 2925
rect 1503 2920 1513 2925
rect 1702 2943 1704 2948
rect 1706 2943 1716 2948
rect 1653 2935 1654 2940
rect 1656 2935 1657 2940
rect 1663 2935 1664 2940
rect 1666 2935 1667 2940
rect 2174 2939 2176 2944
rect 2178 2939 2188 2944
rect 2377 2962 2379 2967
rect 2381 2962 2391 2967
rect 2328 2954 2329 2959
rect 2331 2954 2332 2959
rect 2338 2954 2339 2959
rect 2341 2954 2342 2959
rect 2222 2930 2223 2940
rect 2225 2930 2233 2940
rect 2235 2930 2236 2940
rect 2270 2936 2272 2941
rect 2274 2936 2284 2941
rect 1547 2911 1548 2921
rect 1550 2911 1558 2921
rect 1560 2911 1561 2921
rect 1595 2917 1597 2922
rect 1599 2917 1609 2922
rect 2209 2851 2210 2861
rect 2212 2851 2220 2861
rect 2222 2851 2223 2861
rect 2257 2857 2259 2862
rect 2261 2857 2271 2862
rect 989 2820 990 2830
rect 992 2820 1000 2830
rect 1002 2820 1003 2830
rect 1037 2826 1039 2831
rect 1041 2826 1051 2831
rect 1539 2821 1540 2831
rect 1542 2821 1550 2831
rect 1552 2821 1553 2831
rect 1587 2827 1589 2832
rect 1591 2827 1601 2832
rect 602 2800 603 2810
rect 605 2800 613 2810
rect 615 2800 616 2810
rect 650 2806 652 2811
rect 654 2806 664 2811
<< pdiffusion >>
rect 2522 3884 2523 3894
rect 2525 3884 2527 3894
rect 2531 3884 2533 3894
rect 2535 3884 2536 3894
rect 1900 3866 1901 3876
rect 1903 3866 1905 3876
rect 1909 3866 1911 3876
rect 1913 3866 1914 3876
rect 2476 3874 2478 3884
rect 2480 3874 2490 3884
rect 1854 3856 1856 3866
rect 1858 3856 1868 3866
rect 1179 3840 1180 3850
rect 1182 3840 1184 3850
rect 1188 3840 1190 3850
rect 1192 3840 1193 3850
rect 1133 3830 1135 3840
rect 1137 3830 1147 3840
rect 1227 3837 1229 3847
rect 1231 3837 1241 3847
rect 1948 3863 1950 3873
rect 1952 3863 1962 3873
rect 2570 3881 2572 3891
rect 2574 3881 2584 3891
rect 2008 3820 2009 3840
rect 2011 3820 2019 3840
rect 2021 3820 2022 3840
rect 2630 3838 2631 3858
rect 2633 3838 2641 3858
rect 2643 3838 2644 3858
rect 2679 3841 2681 3851
rect 2683 3841 2693 3851
rect 2057 3823 2059 3833
rect 2061 3823 2071 3833
rect 1287 3794 1288 3814
rect 1290 3794 1298 3814
rect 1300 3794 1301 3814
rect 1336 3797 1338 3807
rect 1340 3797 1350 3807
rect 1854 3800 1856 3810
rect 1858 3800 1868 3810
rect 1902 3800 1903 3810
rect 1905 3800 1907 3810
rect 1911 3800 1913 3810
rect 1915 3800 1916 3810
rect 1133 3774 1135 3784
rect 1137 3774 1147 3784
rect 1181 3774 1182 3784
rect 1184 3774 1186 3784
rect 1190 3774 1192 3784
rect 1194 3774 1195 3784
rect 1229 3771 1231 3781
rect 1233 3771 1243 3781
rect 1950 3797 1952 3807
rect 1954 3797 1964 3807
rect 2476 3818 2478 3828
rect 2480 3818 2490 3828
rect 2524 3818 2525 3828
rect 2527 3818 2529 3828
rect 2533 3818 2535 3828
rect 2537 3818 2538 3828
rect 2572 3815 2574 3825
rect 2576 3815 2586 3825
rect 634 3594 635 3604
rect 637 3594 639 3604
rect 643 3594 645 3604
rect 647 3594 648 3604
rect 588 3584 590 3594
rect 592 3584 602 3594
rect 682 3591 684 3601
rect 686 3591 696 3601
rect 742 3548 743 3568
rect 745 3548 753 3568
rect 755 3548 756 3568
rect 791 3551 793 3561
rect 795 3551 805 3561
rect 588 3528 590 3538
rect 592 3528 602 3538
rect 636 3528 637 3538
rect 639 3528 641 3538
rect 645 3528 647 3538
rect 649 3528 650 3538
rect 684 3525 686 3535
rect 688 3525 698 3535
rect 1974 3488 1975 3498
rect 1977 3488 1979 3498
rect 1983 3488 1985 3498
rect 1987 3488 1988 3498
rect 2022 3485 2024 3495
rect 2026 3485 2036 3495
rect 2113 3429 2114 3449
rect 2116 3429 2124 3449
rect 2126 3429 2127 3449
rect 2162 3432 2164 3442
rect 2166 3432 2176 3442
rect 1973 3365 1974 3375
rect 1976 3365 1978 3375
rect 1982 3365 1984 3375
rect 1986 3365 1987 3375
rect 2021 3362 2023 3372
rect 2025 3362 2035 3372
rect 1489 3332 1490 3342
rect 1492 3332 1494 3342
rect 1498 3332 1500 3342
rect 1502 3332 1503 3342
rect 1537 3329 1539 3339
rect 1541 3329 1551 3339
rect 2289 3309 2290 3329
rect 2292 3309 2300 3329
rect 2302 3309 2303 3329
rect 2338 3312 2340 3322
rect 2342 3312 2352 3322
rect 2474 3318 2475 3338
rect 2477 3318 2485 3338
rect 2487 3318 2488 3338
rect 2523 3321 2525 3331
rect 2527 3321 2537 3331
rect 1621 3284 1622 3304
rect 1624 3284 1632 3304
rect 1634 3284 1635 3304
rect 1670 3287 1672 3297
rect 1674 3287 1684 3297
rect 1737 3245 1738 3265
rect 1740 3245 1748 3265
rect 1750 3245 1751 3265
rect 1786 3248 1788 3258
rect 1790 3248 1800 3258
rect 1488 3226 1489 3236
rect 1491 3226 1493 3236
rect 1497 3226 1499 3236
rect 1501 3226 1502 3236
rect 917 3215 918 3225
rect 920 3215 922 3225
rect 926 3215 928 3225
rect 930 3215 931 3225
rect 965 3212 967 3222
rect 969 3212 979 3222
rect 1536 3223 1538 3233
rect 1540 3223 1550 3233
rect 1978 3242 1979 3252
rect 1981 3242 1983 3252
rect 1987 3242 1989 3252
rect 1991 3242 1992 3252
rect 2026 3239 2028 3249
rect 2030 3239 2040 3249
rect 1625 3182 1626 3202
rect 1628 3182 1636 3202
rect 1638 3182 1639 3202
rect 1674 3185 1676 3195
rect 1678 3185 1688 3195
rect 2112 3185 2113 3205
rect 2115 3185 2123 3205
rect 2125 3185 2126 3205
rect 2161 3188 2163 3198
rect 2165 3188 2175 3198
rect 1043 3141 1044 3161
rect 1046 3141 1054 3161
rect 1056 3141 1057 3161
rect 1092 3144 1094 3154
rect 1096 3144 1106 3154
rect 1158 3151 1159 3171
rect 1161 3151 1169 3171
rect 1171 3151 1172 3171
rect 1207 3154 1209 3164
rect 1211 3154 1221 3164
rect 1492 3129 1493 3139
rect 1495 3129 1497 3139
rect 1501 3129 1503 3139
rect 1505 3129 1506 3139
rect 583 3097 584 3107
rect 586 3097 588 3107
rect 592 3097 594 3107
rect 596 3097 597 3107
rect 631 3094 633 3104
rect 635 3094 645 3104
rect 687 3093 688 3113
rect 690 3093 698 3113
rect 700 3093 701 3113
rect 922 3106 923 3116
rect 925 3106 927 3116
rect 931 3106 933 3116
rect 935 3106 936 3116
rect 736 3096 738 3106
rect 740 3096 750 3106
rect 970 3103 972 3113
rect 974 3103 984 3113
rect 1540 3126 1542 3136
rect 1544 3126 1554 3136
rect 1977 3114 1978 3124
rect 1980 3114 1982 3124
rect 1986 3114 1988 3124
rect 1990 3114 1991 3124
rect 2025 3111 2027 3121
rect 2029 3111 2039 3121
rect 2220 3025 2221 3035
rect 2223 3025 2225 3035
rect 2229 3025 2231 3035
rect 2233 3025 2234 3035
rect 632 3004 633 3014
rect 635 3004 637 3014
rect 641 3004 643 3014
rect 645 3004 646 3014
rect 586 2994 588 3004
rect 590 2994 600 3004
rect 680 3001 682 3011
rect 684 3001 694 3011
rect 984 3006 985 3016
rect 987 3006 989 3016
rect 993 3006 995 3016
rect 997 3006 998 3016
rect 938 2996 940 3006
rect 942 2996 952 3006
rect 1032 3003 1034 3013
rect 1036 3003 1046 3013
rect 1545 3006 1546 3016
rect 1548 3006 1550 3016
rect 1554 3006 1556 3016
rect 1558 3006 1559 3016
rect 2174 3015 2176 3025
rect 2178 3015 2188 3025
rect 1499 2996 1501 3006
rect 1503 2996 1513 3006
rect 740 2958 741 2978
rect 743 2958 751 2978
rect 753 2958 754 2978
rect 1593 3003 1595 3013
rect 1597 3003 1607 3013
rect 2268 3022 2270 3032
rect 2272 3022 2282 3032
rect 789 2961 791 2971
rect 793 2961 803 2971
rect 586 2938 588 2948
rect 590 2938 600 2948
rect 634 2938 635 2948
rect 637 2938 639 2948
rect 643 2938 645 2948
rect 647 2938 648 2948
rect 682 2935 684 2945
rect 686 2935 696 2945
rect 1092 2960 1093 2980
rect 1095 2960 1103 2980
rect 1105 2960 1106 2980
rect 1141 2963 1143 2973
rect 1145 2963 1155 2973
rect 938 2940 940 2950
rect 942 2940 952 2950
rect 986 2940 987 2950
rect 989 2940 991 2950
rect 995 2940 997 2950
rect 999 2940 1000 2950
rect 1034 2937 1036 2947
rect 1038 2937 1048 2947
rect 1653 2960 1654 2980
rect 1656 2960 1664 2980
rect 1666 2960 1667 2980
rect 2328 2979 2329 2999
rect 2331 2979 2339 2999
rect 2341 2979 2342 2999
rect 2377 2982 2379 2992
rect 2381 2982 2391 2992
rect 1702 2963 1704 2973
rect 1706 2963 1716 2973
rect 1499 2940 1501 2950
rect 1503 2940 1513 2950
rect 1547 2940 1548 2950
rect 1550 2940 1552 2950
rect 1556 2940 1558 2950
rect 1560 2940 1561 2950
rect 1595 2937 1597 2947
rect 1599 2937 1609 2947
rect 2174 2959 2176 2969
rect 2178 2959 2188 2969
rect 2222 2959 2223 2969
rect 2225 2959 2227 2969
rect 2231 2959 2233 2969
rect 2235 2959 2236 2969
rect 2270 2956 2272 2966
rect 2274 2956 2284 2966
rect 2209 2880 2210 2890
rect 2212 2880 2214 2890
rect 2218 2880 2220 2890
rect 2222 2880 2223 2890
rect 2257 2877 2259 2887
rect 2261 2877 2271 2887
rect 989 2849 990 2859
rect 992 2849 994 2859
rect 998 2849 1000 2859
rect 1002 2849 1003 2859
rect 602 2829 603 2839
rect 605 2829 607 2839
rect 611 2829 613 2839
rect 615 2829 616 2839
rect 650 2826 652 2836
rect 654 2826 664 2836
rect 1037 2846 1039 2856
rect 1041 2846 1051 2856
rect 1539 2850 1540 2860
rect 1542 2850 1544 2860
rect 1548 2850 1550 2860
rect 1552 2850 1553 2860
rect 1587 2847 1589 2857
rect 1591 2847 1601 2857
<< ndcontact >>
rect 2472 3854 2476 3859
rect 2490 3854 2494 3859
rect 2518 3855 2522 3865
rect 2536 3855 2540 3865
rect 2566 3861 2570 3866
rect 2584 3861 2588 3866
rect 1850 3836 1854 3841
rect 1868 3836 1872 3841
rect 1896 3837 1900 3847
rect 1914 3837 1918 3847
rect 1944 3843 1948 3848
rect 1962 3843 1966 3848
rect 1129 3810 1133 3815
rect 1147 3810 1151 3815
rect 1175 3811 1179 3821
rect 1193 3811 1197 3821
rect 1223 3817 1227 3822
rect 1241 3817 1245 3822
rect 1129 3754 1133 3759
rect 1147 3754 1151 3759
rect 1332 3777 1336 3782
rect 1350 3777 1354 3782
rect 1850 3780 1854 3785
rect 1868 3780 1872 3785
rect 2053 3803 2057 3808
rect 2071 3803 2075 3808
rect 2004 3795 2008 3800
rect 2012 3795 2018 3800
rect 2022 3795 2026 3800
rect 2472 3798 2476 3803
rect 2490 3798 2494 3803
rect 2675 3821 2679 3826
rect 2693 3821 2697 3826
rect 2626 3813 2630 3818
rect 2634 3813 2640 3818
rect 2644 3813 2648 3818
rect 2520 3789 2524 3799
rect 2538 3789 2542 3799
rect 2568 3795 2572 3800
rect 2586 3795 2590 3800
rect 1283 3769 1287 3774
rect 1291 3769 1297 3774
rect 1301 3769 1305 3774
rect 1898 3771 1902 3781
rect 1916 3771 1920 3781
rect 1946 3777 1950 3782
rect 1964 3777 1968 3782
rect 1177 3745 1181 3755
rect 1195 3745 1199 3755
rect 1225 3751 1229 3756
rect 1243 3751 1247 3756
rect 584 3564 588 3569
rect 602 3564 606 3569
rect 630 3565 634 3575
rect 648 3565 652 3575
rect 678 3571 682 3576
rect 696 3571 700 3576
rect 584 3508 588 3513
rect 602 3508 606 3513
rect 787 3531 791 3536
rect 805 3531 809 3536
rect 738 3523 742 3528
rect 746 3523 752 3528
rect 756 3523 760 3528
rect 632 3499 636 3509
rect 650 3499 654 3509
rect 680 3505 684 3510
rect 698 3505 702 3510
rect 1970 3459 1974 3469
rect 1988 3459 1992 3469
rect 2018 3465 2022 3470
rect 2036 3465 2040 3470
rect 2158 3412 2162 3417
rect 2176 3412 2180 3417
rect 2109 3404 2113 3409
rect 2117 3404 2123 3409
rect 2127 3404 2131 3409
rect 1969 3336 1973 3346
rect 1987 3336 1991 3346
rect 2017 3342 2021 3347
rect 2035 3342 2039 3347
rect 1485 3303 1489 3313
rect 1503 3303 1507 3313
rect 1533 3309 1537 3314
rect 1551 3309 1555 3314
rect 2519 3301 2523 3306
rect 2537 3301 2541 3306
rect 2334 3292 2338 3297
rect 2352 3292 2356 3297
rect 2470 3293 2474 3298
rect 2478 3293 2484 3298
rect 2488 3293 2492 3298
rect 2285 3284 2289 3289
rect 2293 3284 2299 3289
rect 2303 3284 2307 3289
rect 1666 3267 1670 3272
rect 1684 3267 1688 3272
rect 1617 3259 1621 3264
rect 1625 3259 1631 3264
rect 1635 3259 1639 3264
rect 1782 3228 1786 3233
rect 1800 3228 1804 3233
rect 1733 3220 1737 3225
rect 1741 3220 1747 3225
rect 1751 3220 1755 3225
rect 1974 3213 1978 3223
rect 1992 3213 1996 3223
rect 2022 3219 2026 3224
rect 2040 3219 2044 3224
rect 1484 3197 1488 3207
rect 1502 3197 1506 3207
rect 1532 3203 1536 3208
rect 1550 3203 1554 3208
rect 913 3186 917 3196
rect 931 3186 935 3196
rect 961 3192 965 3197
rect 979 3192 983 3197
rect 1670 3165 1674 3170
rect 1688 3165 1692 3170
rect 2157 3168 2161 3173
rect 2175 3168 2179 3173
rect 1621 3157 1625 3162
rect 1629 3157 1635 3162
rect 1639 3157 1643 3162
rect 2108 3160 2112 3165
rect 2116 3160 2122 3165
rect 2126 3160 2130 3165
rect 1203 3134 1207 3139
rect 1221 3134 1225 3139
rect 1088 3124 1092 3129
rect 1106 3124 1110 3129
rect 1154 3126 1158 3131
rect 1162 3126 1168 3131
rect 1172 3126 1176 3131
rect 1039 3116 1043 3121
rect 1047 3116 1053 3121
rect 1057 3116 1061 3121
rect 579 3068 583 3078
rect 597 3068 601 3078
rect 627 3074 631 3079
rect 645 3074 649 3079
rect 1488 3100 1492 3110
rect 1506 3100 1510 3110
rect 1536 3106 1540 3111
rect 1554 3106 1558 3111
rect 732 3076 736 3081
rect 750 3076 754 3081
rect 918 3077 922 3087
rect 936 3077 940 3087
rect 966 3083 970 3088
rect 984 3083 988 3088
rect 1973 3085 1977 3095
rect 1991 3085 1995 3095
rect 2021 3091 2025 3096
rect 2039 3091 2043 3096
rect 683 3068 687 3073
rect 691 3068 697 3073
rect 701 3068 705 3073
rect 582 2974 586 2979
rect 600 2974 604 2979
rect 628 2975 632 2985
rect 646 2975 650 2985
rect 676 2981 680 2986
rect 694 2981 698 2986
rect 934 2976 938 2981
rect 952 2976 956 2981
rect 980 2977 984 2987
rect 998 2977 1002 2987
rect 1028 2983 1032 2988
rect 1046 2983 1050 2988
rect 2170 2995 2174 3000
rect 2188 2995 2192 3000
rect 2216 2996 2220 3006
rect 2234 2996 2238 3006
rect 2264 3002 2268 3007
rect 2282 3002 2286 3007
rect 582 2918 586 2923
rect 600 2918 604 2923
rect 1495 2976 1499 2981
rect 1513 2976 1517 2981
rect 1541 2977 1545 2987
rect 1559 2977 1563 2987
rect 1589 2983 1593 2988
rect 1607 2983 1611 2988
rect 785 2941 789 2946
rect 803 2941 807 2946
rect 736 2933 740 2938
rect 744 2933 750 2938
rect 754 2933 758 2938
rect 934 2920 938 2925
rect 952 2920 956 2925
rect 1137 2943 1141 2948
rect 1155 2943 1159 2948
rect 1088 2935 1092 2940
rect 1096 2935 1102 2940
rect 1106 2935 1110 2940
rect 630 2909 634 2919
rect 648 2909 652 2919
rect 678 2915 682 2920
rect 696 2915 700 2920
rect 982 2911 986 2921
rect 1000 2911 1004 2921
rect 1030 2917 1034 2922
rect 1048 2917 1052 2922
rect 1495 2920 1499 2925
rect 1513 2920 1517 2925
rect 1698 2943 1702 2948
rect 1716 2943 1720 2948
rect 1649 2935 1653 2940
rect 1657 2935 1663 2940
rect 1667 2935 1671 2940
rect 2170 2939 2174 2944
rect 2188 2939 2192 2944
rect 2373 2962 2377 2967
rect 2391 2962 2395 2967
rect 2324 2954 2328 2959
rect 2332 2954 2338 2959
rect 2342 2954 2346 2959
rect 2218 2930 2222 2940
rect 2236 2930 2240 2940
rect 2266 2936 2270 2941
rect 2284 2936 2288 2941
rect 1543 2911 1547 2921
rect 1561 2911 1565 2921
rect 1591 2917 1595 2922
rect 1609 2917 1613 2922
rect 2205 2851 2209 2861
rect 2223 2851 2227 2861
rect 2253 2857 2257 2862
rect 2271 2857 2275 2862
rect 985 2820 989 2830
rect 1003 2820 1007 2830
rect 1033 2826 1037 2831
rect 1051 2826 1055 2831
rect 1535 2821 1539 2831
rect 1553 2821 1557 2831
rect 1583 2827 1587 2832
rect 1601 2827 1605 2832
rect 598 2800 602 2810
rect 616 2800 620 2810
rect 646 2806 650 2811
rect 664 2806 668 2811
<< pdcontact >>
rect 2518 3884 2522 3894
rect 2527 3884 2531 3894
rect 2536 3884 2540 3894
rect 1896 3866 1900 3876
rect 1905 3866 1909 3876
rect 1914 3866 1918 3876
rect 2472 3874 2476 3884
rect 2490 3874 2494 3884
rect 1850 3856 1854 3866
rect 1868 3856 1872 3866
rect 1175 3840 1179 3850
rect 1184 3840 1188 3850
rect 1193 3840 1197 3850
rect 1129 3830 1133 3840
rect 1147 3830 1151 3840
rect 1223 3837 1227 3847
rect 1241 3837 1245 3847
rect 1944 3863 1948 3873
rect 1962 3863 1966 3873
rect 2566 3881 2570 3891
rect 2584 3881 2588 3891
rect 2004 3820 2008 3840
rect 2022 3820 2026 3840
rect 2626 3838 2630 3858
rect 2644 3838 2648 3858
rect 2675 3841 2679 3851
rect 2693 3841 2697 3851
rect 2053 3823 2057 3833
rect 2071 3823 2075 3833
rect 1283 3794 1287 3814
rect 1301 3794 1305 3814
rect 1332 3797 1336 3807
rect 1350 3797 1354 3807
rect 1850 3800 1854 3810
rect 1868 3800 1872 3810
rect 1898 3800 1902 3810
rect 1907 3800 1911 3810
rect 1916 3800 1920 3810
rect 1129 3774 1133 3784
rect 1147 3774 1151 3784
rect 1177 3774 1181 3784
rect 1186 3774 1190 3784
rect 1195 3774 1199 3784
rect 1225 3771 1229 3781
rect 1243 3771 1247 3781
rect 1946 3797 1950 3807
rect 1964 3797 1968 3807
rect 2472 3818 2476 3828
rect 2490 3818 2494 3828
rect 2520 3818 2524 3828
rect 2529 3818 2533 3828
rect 2538 3818 2542 3828
rect 2568 3815 2572 3825
rect 2586 3815 2590 3825
rect 630 3594 634 3604
rect 639 3594 643 3604
rect 648 3594 652 3604
rect 584 3584 588 3594
rect 602 3584 606 3594
rect 678 3591 682 3601
rect 696 3591 700 3601
rect 738 3548 742 3568
rect 756 3548 760 3568
rect 787 3551 791 3561
rect 805 3551 809 3561
rect 584 3528 588 3538
rect 602 3528 606 3538
rect 632 3528 636 3538
rect 641 3528 645 3538
rect 650 3528 654 3538
rect 680 3525 684 3535
rect 698 3525 702 3535
rect 1970 3488 1974 3498
rect 1979 3488 1983 3498
rect 1988 3488 1992 3498
rect 2018 3485 2022 3495
rect 2036 3485 2040 3495
rect 2109 3429 2113 3449
rect 2127 3429 2131 3449
rect 2158 3432 2162 3442
rect 2176 3432 2180 3442
rect 1969 3365 1973 3375
rect 1978 3365 1982 3375
rect 1987 3365 1991 3375
rect 2017 3362 2021 3372
rect 2035 3362 2039 3372
rect 1485 3332 1489 3342
rect 1494 3332 1498 3342
rect 1503 3332 1507 3342
rect 1533 3329 1537 3339
rect 1551 3329 1555 3339
rect 2285 3309 2289 3329
rect 2303 3309 2307 3329
rect 2334 3312 2338 3322
rect 2352 3312 2356 3322
rect 2470 3318 2474 3338
rect 2488 3318 2492 3338
rect 2519 3321 2523 3331
rect 2537 3321 2541 3331
rect 1617 3284 1621 3304
rect 1635 3284 1639 3304
rect 1666 3287 1670 3297
rect 1684 3287 1688 3297
rect 1733 3245 1737 3265
rect 1751 3245 1755 3265
rect 1782 3248 1786 3258
rect 1800 3248 1804 3258
rect 1484 3226 1488 3236
rect 1493 3226 1497 3236
rect 1502 3226 1506 3236
rect 913 3215 917 3225
rect 922 3215 926 3225
rect 931 3215 935 3225
rect 961 3212 965 3222
rect 979 3212 983 3222
rect 1532 3223 1536 3233
rect 1550 3223 1554 3233
rect 1974 3242 1978 3252
rect 1983 3242 1987 3252
rect 1992 3242 1996 3252
rect 2022 3239 2026 3249
rect 2040 3239 2044 3249
rect 1621 3182 1625 3202
rect 1639 3182 1643 3202
rect 1670 3185 1674 3195
rect 1688 3185 1692 3195
rect 2108 3185 2112 3205
rect 2126 3185 2130 3205
rect 2157 3188 2161 3198
rect 2175 3188 2179 3198
rect 1039 3141 1043 3161
rect 1057 3141 1061 3161
rect 1088 3144 1092 3154
rect 1106 3144 1110 3154
rect 1154 3151 1158 3171
rect 1172 3151 1176 3171
rect 1203 3154 1207 3164
rect 1221 3154 1225 3164
rect 1488 3129 1492 3139
rect 1497 3129 1501 3139
rect 1506 3129 1510 3139
rect 579 3097 583 3107
rect 588 3097 592 3107
rect 597 3097 601 3107
rect 627 3094 631 3104
rect 645 3094 649 3104
rect 683 3093 687 3113
rect 701 3093 705 3113
rect 918 3106 922 3116
rect 927 3106 931 3116
rect 936 3106 940 3116
rect 732 3096 736 3106
rect 750 3096 754 3106
rect 966 3103 970 3113
rect 984 3103 988 3113
rect 1536 3126 1540 3136
rect 1554 3126 1558 3136
rect 1973 3114 1977 3124
rect 1982 3114 1986 3124
rect 1991 3114 1995 3124
rect 2021 3111 2025 3121
rect 2039 3111 2043 3121
rect 2216 3025 2220 3035
rect 2225 3025 2229 3035
rect 2234 3025 2238 3035
rect 628 3004 632 3014
rect 637 3004 641 3014
rect 646 3004 650 3014
rect 582 2994 586 3004
rect 600 2994 604 3004
rect 676 3001 680 3011
rect 694 3001 698 3011
rect 980 3006 984 3016
rect 989 3006 993 3016
rect 998 3006 1002 3016
rect 934 2996 938 3006
rect 952 2996 956 3006
rect 1028 3003 1032 3013
rect 1046 3003 1050 3013
rect 1541 3006 1545 3016
rect 1550 3006 1554 3016
rect 1559 3006 1563 3016
rect 2170 3015 2174 3025
rect 2188 3015 2192 3025
rect 1495 2996 1499 3006
rect 1513 2996 1517 3006
rect 736 2958 740 2978
rect 754 2958 758 2978
rect 1589 3003 1593 3013
rect 1607 3003 1611 3013
rect 2264 3022 2268 3032
rect 2282 3022 2286 3032
rect 785 2961 789 2971
rect 803 2961 807 2971
rect 582 2938 586 2948
rect 600 2938 604 2948
rect 630 2938 634 2948
rect 639 2938 643 2948
rect 648 2938 652 2948
rect 678 2935 682 2945
rect 696 2935 700 2945
rect 1088 2960 1092 2980
rect 1106 2960 1110 2980
rect 1137 2963 1141 2973
rect 1155 2963 1159 2973
rect 934 2940 938 2950
rect 952 2940 956 2950
rect 982 2940 986 2950
rect 991 2940 995 2950
rect 1000 2940 1004 2950
rect 1030 2937 1034 2947
rect 1048 2937 1052 2947
rect 1649 2960 1653 2980
rect 1667 2960 1671 2980
rect 2324 2979 2328 2999
rect 2342 2979 2346 2999
rect 2373 2982 2377 2992
rect 2391 2982 2395 2992
rect 1698 2963 1702 2973
rect 1716 2963 1720 2973
rect 1495 2940 1499 2950
rect 1513 2940 1517 2950
rect 1543 2940 1547 2950
rect 1552 2940 1556 2950
rect 1561 2940 1565 2950
rect 1591 2937 1595 2947
rect 1609 2937 1613 2947
rect 2170 2959 2174 2969
rect 2188 2959 2192 2969
rect 2218 2959 2222 2969
rect 2227 2959 2231 2969
rect 2236 2959 2240 2969
rect 2266 2956 2270 2966
rect 2284 2956 2288 2966
rect 2205 2880 2209 2890
rect 2214 2880 2218 2890
rect 2223 2880 2227 2890
rect 2253 2877 2257 2887
rect 2271 2877 2275 2887
rect 985 2849 989 2859
rect 994 2849 998 2859
rect 1003 2849 1007 2859
rect 598 2829 602 2839
rect 607 2829 611 2839
rect 616 2829 620 2839
rect 646 2826 650 2836
rect 664 2826 668 2836
rect 1033 2846 1037 2856
rect 1051 2846 1055 2856
rect 1535 2850 1539 2860
rect 1544 2850 1548 2860
rect 1553 2850 1557 2860
rect 1583 2847 1587 2857
rect 1601 2847 1605 2857
<< polysilicon >>
rect 2523 3894 2525 3897
rect 2533 3894 2535 3897
rect 2478 3884 2480 3887
rect 2572 3891 2574 3894
rect 1901 3876 1903 3879
rect 1911 3876 1913 3879
rect 1856 3866 1858 3869
rect 1950 3873 1952 3876
rect 1180 3850 1182 3853
rect 1190 3850 1192 3853
rect 1135 3840 1137 3843
rect 1229 3847 1231 3850
rect 1135 3815 1137 3830
rect 1180 3821 1182 3840
rect 1190 3821 1192 3840
rect 1856 3841 1858 3856
rect 1901 3847 1903 3866
rect 1911 3847 1913 3866
rect 1950 3848 1952 3863
rect 2478 3859 2480 3874
rect 2523 3865 2525 3884
rect 2533 3865 2535 3884
rect 2572 3866 2574 3881
rect 2572 3858 2574 3861
rect 2631 3858 2633 3861
rect 2641 3858 2643 3861
rect 2478 3851 2480 3854
rect 2523 3852 2525 3855
rect 2533 3852 2535 3855
rect 1229 3822 1231 3837
rect 1950 3840 1952 3843
rect 2009 3840 2011 3843
rect 2019 3840 2021 3843
rect 1856 3833 1858 3836
rect 1901 3834 1903 3837
rect 1911 3834 1913 3837
rect 2681 3851 2683 3854
rect 2059 3833 2061 3836
rect 2478 3828 2480 3831
rect 2525 3828 2527 3831
rect 2535 3828 2537 3831
rect 1229 3814 1231 3817
rect 1288 3814 1290 3817
rect 1298 3814 1300 3817
rect 1135 3807 1137 3810
rect 1180 3808 1182 3811
rect 1190 3808 1192 3811
rect 1856 3810 1858 3813
rect 1903 3810 1905 3813
rect 1913 3810 1915 3813
rect 1338 3807 1340 3810
rect 1952 3807 1954 3810
rect 1135 3784 1137 3787
rect 1182 3784 1184 3787
rect 1192 3784 1194 3787
rect 1231 3781 1233 3784
rect 1135 3759 1137 3774
rect 1182 3755 1184 3774
rect 1192 3755 1194 3774
rect 1288 3774 1290 3794
rect 1298 3774 1300 3794
rect 1338 3782 1340 3797
rect 1856 3785 1858 3800
rect 1903 3781 1905 3800
rect 1913 3781 1915 3800
rect 2009 3800 2011 3820
rect 2019 3800 2021 3820
rect 2059 3808 2061 3823
rect 2574 3825 2576 3828
rect 2478 3803 2480 3818
rect 2059 3800 2061 3803
rect 1952 3782 1954 3797
rect 2525 3799 2527 3818
rect 2535 3799 2537 3818
rect 2631 3818 2633 3838
rect 2641 3818 2643 3838
rect 2681 3826 2683 3841
rect 2681 3818 2683 3821
rect 2574 3800 2576 3815
rect 2631 3810 2633 3813
rect 2641 3810 2643 3813
rect 2478 3795 2480 3798
rect 2009 3792 2011 3795
rect 2019 3792 2021 3795
rect 2574 3792 2576 3795
rect 2525 3786 2527 3789
rect 2535 3786 2537 3789
rect 1856 3777 1858 3780
rect 1338 3774 1340 3777
rect 1231 3756 1233 3771
rect 1952 3774 1954 3777
rect 1288 3766 1290 3769
rect 1298 3766 1300 3769
rect 1903 3768 1905 3771
rect 1913 3768 1915 3771
rect 1135 3751 1137 3754
rect 1231 3748 1233 3751
rect 1182 3742 1184 3745
rect 1192 3742 1194 3745
rect 635 3604 637 3607
rect 645 3604 647 3607
rect 590 3594 592 3597
rect 684 3601 686 3604
rect 590 3569 592 3584
rect 635 3575 637 3594
rect 645 3575 647 3594
rect 684 3576 686 3591
rect 684 3568 686 3571
rect 743 3568 745 3571
rect 753 3568 755 3571
rect 590 3561 592 3564
rect 635 3562 637 3565
rect 645 3562 647 3565
rect 793 3561 795 3564
rect 590 3538 592 3541
rect 637 3538 639 3541
rect 647 3538 649 3541
rect 686 3535 688 3538
rect 590 3513 592 3528
rect 637 3509 639 3528
rect 647 3509 649 3528
rect 743 3528 745 3548
rect 753 3528 755 3548
rect 793 3536 795 3551
rect 793 3528 795 3531
rect 686 3510 688 3525
rect 743 3520 745 3523
rect 753 3520 755 3523
rect 590 3505 592 3508
rect 686 3502 688 3505
rect 637 3496 639 3499
rect 647 3496 649 3499
rect 1975 3498 1977 3501
rect 1985 3498 1987 3501
rect 2024 3495 2026 3498
rect 1975 3469 1977 3488
rect 1985 3469 1987 3488
rect 2024 3470 2026 3485
rect 2024 3462 2026 3465
rect 1975 3456 1977 3459
rect 1985 3456 1987 3459
rect 2114 3449 2116 3452
rect 2124 3449 2126 3452
rect 2164 3442 2166 3445
rect 2114 3409 2116 3429
rect 2124 3409 2126 3429
rect 2164 3417 2166 3432
rect 2164 3409 2166 3412
rect 2114 3401 2116 3404
rect 2124 3401 2126 3404
rect 1974 3375 1976 3378
rect 1984 3375 1986 3378
rect 2023 3372 2025 3375
rect 1974 3346 1976 3365
rect 1984 3346 1986 3365
rect 2023 3347 2025 3362
rect 1490 3342 1492 3345
rect 1500 3342 1502 3345
rect 1539 3339 1541 3342
rect 1490 3313 1492 3332
rect 1500 3313 1502 3332
rect 2023 3339 2025 3342
rect 2475 3338 2477 3341
rect 2485 3338 2487 3341
rect 1974 3333 1976 3336
rect 1984 3333 1986 3336
rect 2290 3329 2292 3332
rect 2300 3329 2302 3332
rect 1539 3314 1541 3329
rect 2340 3322 2342 3325
rect 2525 3331 2527 3334
rect 1539 3306 1541 3309
rect 1622 3304 1624 3307
rect 1632 3304 1634 3307
rect 1490 3300 1492 3303
rect 1500 3300 1502 3303
rect 1672 3297 1674 3300
rect 2290 3289 2292 3309
rect 2300 3289 2302 3309
rect 2340 3297 2342 3312
rect 2475 3298 2477 3318
rect 2485 3298 2487 3318
rect 2525 3306 2527 3321
rect 2525 3298 2527 3301
rect 2340 3289 2342 3292
rect 2475 3290 2477 3293
rect 2485 3290 2487 3293
rect 1622 3264 1624 3284
rect 1632 3264 1634 3284
rect 1672 3272 1674 3287
rect 2290 3281 2292 3284
rect 2300 3281 2302 3284
rect 1672 3264 1674 3267
rect 1738 3265 1740 3268
rect 1748 3265 1750 3268
rect 1622 3256 1624 3259
rect 1632 3256 1634 3259
rect 1788 3258 1790 3261
rect 1979 3252 1981 3255
rect 1989 3252 1991 3255
rect 1489 3236 1491 3239
rect 1499 3236 1501 3239
rect 918 3225 920 3228
rect 928 3225 930 3228
rect 1538 3233 1540 3236
rect 967 3222 969 3225
rect 918 3196 920 3215
rect 928 3196 930 3215
rect 967 3197 969 3212
rect 1489 3207 1491 3226
rect 1499 3207 1501 3226
rect 1738 3225 1740 3245
rect 1748 3225 1750 3245
rect 1788 3233 1790 3248
rect 2028 3249 2030 3252
rect 1788 3225 1790 3228
rect 1538 3208 1540 3223
rect 1979 3223 1981 3242
rect 1989 3223 1991 3242
rect 2028 3224 2030 3239
rect 1738 3217 1740 3220
rect 1748 3217 1750 3220
rect 2028 3216 2030 3219
rect 1979 3210 1981 3213
rect 1989 3210 1991 3213
rect 2113 3205 2115 3208
rect 2123 3205 2125 3208
rect 1538 3200 1540 3203
rect 1626 3202 1628 3205
rect 1636 3202 1638 3205
rect 1489 3194 1491 3197
rect 1499 3194 1501 3197
rect 967 3189 969 3192
rect 918 3183 920 3186
rect 928 3183 930 3186
rect 1676 3195 1678 3198
rect 2163 3198 2165 3201
rect 1159 3171 1161 3174
rect 1169 3171 1171 3174
rect 1044 3161 1046 3164
rect 1054 3161 1056 3164
rect 1094 3154 1096 3157
rect 1209 3164 1211 3167
rect 1626 3162 1628 3182
rect 1636 3162 1638 3182
rect 1676 3170 1678 3185
rect 2113 3165 2115 3185
rect 2123 3165 2125 3185
rect 2163 3173 2165 3188
rect 2163 3165 2165 3168
rect 1676 3162 1678 3165
rect 2113 3157 2115 3160
rect 2123 3157 2125 3160
rect 1626 3154 1628 3157
rect 1636 3154 1638 3157
rect 1044 3121 1046 3141
rect 1054 3121 1056 3141
rect 1094 3129 1096 3144
rect 1159 3131 1161 3151
rect 1169 3131 1171 3151
rect 1209 3139 1211 3154
rect 1493 3139 1495 3142
rect 1503 3139 1505 3142
rect 1209 3131 1211 3134
rect 1542 3136 1544 3139
rect 1094 3121 1096 3124
rect 1159 3123 1161 3126
rect 1169 3123 1171 3126
rect 923 3116 925 3119
rect 933 3116 935 3119
rect 688 3113 690 3116
rect 698 3113 700 3116
rect 584 3107 586 3110
rect 594 3107 596 3110
rect 633 3104 635 3107
rect 584 3078 586 3097
rect 594 3078 596 3097
rect 633 3079 635 3094
rect 738 3106 740 3109
rect 972 3113 974 3116
rect 1044 3113 1046 3116
rect 1054 3113 1056 3116
rect 633 3071 635 3074
rect 688 3073 690 3093
rect 698 3073 700 3093
rect 738 3081 740 3096
rect 923 3087 925 3106
rect 933 3087 935 3106
rect 1493 3110 1495 3129
rect 1503 3110 1505 3129
rect 1542 3111 1544 3126
rect 1978 3124 1980 3127
rect 1988 3124 1990 3127
rect 2027 3121 2029 3124
rect 972 3088 974 3103
rect 1542 3103 1544 3106
rect 1493 3097 1495 3100
rect 1503 3097 1505 3100
rect 1978 3095 1980 3114
rect 1988 3095 1990 3114
rect 2027 3096 2029 3111
rect 2027 3088 2029 3091
rect 972 3080 974 3083
rect 1978 3082 1980 3085
rect 1988 3082 1990 3085
rect 738 3073 740 3076
rect 923 3074 925 3077
rect 933 3074 935 3077
rect 584 3065 586 3068
rect 594 3065 596 3068
rect 688 3065 690 3068
rect 698 3065 700 3068
rect 2221 3035 2223 3038
rect 2231 3035 2233 3038
rect 2176 3025 2178 3028
rect 2270 3032 2272 3035
rect 633 3014 635 3017
rect 643 3014 645 3017
rect 985 3016 987 3019
rect 995 3016 997 3019
rect 1546 3016 1548 3019
rect 1556 3016 1558 3019
rect 588 3004 590 3007
rect 682 3011 684 3014
rect 588 2979 590 2994
rect 633 2985 635 3004
rect 643 2985 645 3004
rect 940 3006 942 3009
rect 1034 3013 1036 3016
rect 682 2986 684 3001
rect 940 2981 942 2996
rect 985 2987 987 3006
rect 995 2987 997 3006
rect 1501 3006 1503 3009
rect 1595 3013 1597 3016
rect 1034 2988 1036 3003
rect 682 2978 684 2981
rect 741 2978 743 2981
rect 751 2978 753 2981
rect 588 2971 590 2974
rect 633 2972 635 2975
rect 643 2972 645 2975
rect 1034 2980 1036 2983
rect 1093 2980 1095 2983
rect 1103 2980 1105 2983
rect 1501 2981 1503 2996
rect 1546 2987 1548 3006
rect 1556 2987 1558 3006
rect 1595 2988 1597 3003
rect 2176 3000 2178 3015
rect 2221 3006 2223 3025
rect 2231 3006 2233 3025
rect 2270 3007 2272 3022
rect 2270 2999 2272 3002
rect 2329 2999 2331 3002
rect 2339 2999 2341 3002
rect 2176 2992 2178 2995
rect 2221 2993 2223 2996
rect 2231 2993 2233 2996
rect 791 2971 793 2974
rect 940 2973 942 2976
rect 985 2974 987 2977
rect 995 2974 997 2977
rect 588 2948 590 2951
rect 635 2948 637 2951
rect 645 2948 647 2951
rect 684 2945 686 2948
rect 588 2923 590 2938
rect 635 2919 637 2938
rect 645 2919 647 2938
rect 741 2938 743 2958
rect 751 2938 753 2958
rect 791 2946 793 2961
rect 1595 2980 1597 2983
rect 1654 2980 1656 2983
rect 1664 2980 1666 2983
rect 1143 2973 1145 2976
rect 1501 2973 1503 2976
rect 1546 2974 1548 2977
rect 1556 2974 1558 2977
rect 940 2950 942 2953
rect 987 2950 989 2953
rect 997 2950 999 2953
rect 791 2938 793 2941
rect 1036 2947 1038 2950
rect 684 2920 686 2935
rect 741 2930 743 2933
rect 751 2930 753 2933
rect 940 2925 942 2940
rect 987 2921 989 2940
rect 997 2921 999 2940
rect 1093 2940 1095 2960
rect 1103 2940 1105 2960
rect 1143 2948 1145 2963
rect 2379 2992 2381 2995
rect 1704 2973 1706 2976
rect 2176 2969 2178 2972
rect 2223 2969 2225 2972
rect 2233 2969 2235 2972
rect 1501 2950 1503 2953
rect 1548 2950 1550 2953
rect 1558 2950 1560 2953
rect 1143 2940 1145 2943
rect 1597 2947 1599 2950
rect 1036 2922 1038 2937
rect 1093 2932 1095 2935
rect 1103 2932 1105 2935
rect 1501 2925 1503 2940
rect 588 2915 590 2918
rect 940 2917 942 2920
rect 684 2912 686 2915
rect 1548 2921 1550 2940
rect 1558 2921 1560 2940
rect 1654 2940 1656 2960
rect 1664 2940 1666 2960
rect 1704 2948 1706 2963
rect 2272 2966 2274 2969
rect 2176 2944 2178 2959
rect 1704 2940 1706 2943
rect 1597 2922 1599 2937
rect 2223 2940 2225 2959
rect 2233 2940 2235 2959
rect 2329 2959 2331 2979
rect 2339 2959 2341 2979
rect 2379 2967 2381 2982
rect 2379 2959 2381 2962
rect 2272 2941 2274 2956
rect 2329 2951 2331 2954
rect 2339 2951 2341 2954
rect 2176 2936 2178 2939
rect 1654 2932 1656 2935
rect 1664 2932 1666 2935
rect 2272 2933 2274 2936
rect 2223 2927 2225 2930
rect 2233 2927 2235 2930
rect 1501 2917 1503 2920
rect 1036 2914 1038 2917
rect 1597 2914 1599 2917
rect 635 2906 637 2909
rect 645 2906 647 2909
rect 987 2908 989 2911
rect 997 2908 999 2911
rect 1548 2908 1550 2911
rect 1558 2908 1560 2911
rect 2210 2890 2212 2893
rect 2220 2890 2222 2893
rect 2259 2887 2261 2890
rect 990 2859 992 2862
rect 1000 2859 1002 2862
rect 1540 2860 1542 2863
rect 1550 2860 1552 2863
rect 2210 2861 2212 2880
rect 2220 2861 2222 2880
rect 2259 2862 2261 2877
rect 1039 2856 1041 2859
rect 603 2839 605 2842
rect 613 2839 615 2842
rect 652 2836 654 2839
rect 603 2810 605 2829
rect 613 2810 615 2829
rect 990 2830 992 2849
rect 1000 2830 1002 2849
rect 1589 2857 1591 2860
rect 1039 2831 1041 2846
rect 1540 2831 1542 2850
rect 1550 2831 1552 2850
rect 2259 2854 2261 2857
rect 2210 2848 2212 2851
rect 2220 2848 2222 2851
rect 1589 2832 1591 2847
rect 652 2811 654 2826
rect 1039 2823 1041 2826
rect 1589 2824 1591 2827
rect 990 2817 992 2820
rect 1000 2817 1002 2820
rect 1540 2818 1542 2821
rect 1550 2818 1552 2821
rect 652 2803 654 2806
rect 603 2797 605 2800
rect 613 2797 615 2800
<< polycontact >>
rect 1131 3818 1135 3822
rect 1176 3829 1180 3833
rect 1852 3844 1856 3848
rect 1897 3855 1901 3859
rect 1913 3855 1917 3859
rect 1946 3851 1950 3855
rect 2474 3862 2478 3866
rect 2519 3873 2523 3877
rect 2535 3873 2539 3877
rect 2568 3869 2572 3873
rect 1192 3829 1196 3833
rect 1225 3825 1229 3829
rect 2005 3809 2009 3813
rect 1284 3783 1288 3787
rect 1131 3762 1135 3766
rect 1178 3763 1182 3767
rect 1294 3783 1298 3787
rect 1334 3785 1338 3789
rect 1852 3788 1856 3792
rect 1899 3789 1903 3793
rect 2015 3809 2019 3813
rect 2055 3811 2059 3815
rect 2627 3827 2631 3831
rect 2474 3806 2478 3810
rect 2521 3807 2525 3811
rect 1915 3789 1919 3793
rect 1948 3785 1952 3789
rect 2637 3827 2641 3831
rect 2677 3829 2681 3833
rect 2537 3807 2541 3811
rect 2570 3803 2574 3807
rect 1194 3763 1198 3767
rect 1227 3759 1231 3763
rect 586 3572 590 3576
rect 631 3583 635 3587
rect 647 3583 651 3587
rect 680 3579 684 3583
rect 739 3537 743 3541
rect 586 3516 590 3520
rect 633 3517 637 3521
rect 749 3537 753 3541
rect 789 3539 793 3543
rect 649 3517 653 3521
rect 682 3513 686 3517
rect 1971 3476 1975 3481
rect 1987 3477 1991 3481
rect 2020 3473 2024 3477
rect 2110 3418 2114 3422
rect 2120 3418 2124 3422
rect 2160 3420 2164 3424
rect 1970 3354 1974 3358
rect 1986 3354 1990 3358
rect 2019 3350 2023 3354
rect 1486 3321 1490 3325
rect 1502 3321 1506 3325
rect 1535 3317 1539 3321
rect 2286 3298 2290 3302
rect 2296 3298 2300 3302
rect 2336 3300 2340 3304
rect 2471 3307 2475 3311
rect 2481 3307 2485 3311
rect 2521 3309 2525 3313
rect 1618 3273 1622 3277
rect 1628 3273 1632 3277
rect 1668 3275 1672 3279
rect 1734 3234 1738 3238
rect 914 3203 918 3208
rect 1485 3215 1489 3219
rect 930 3204 934 3208
rect 963 3200 967 3204
rect 1744 3234 1748 3238
rect 1784 3236 1788 3240
rect 1975 3231 1979 3235
rect 1501 3215 1505 3219
rect 1534 3211 1538 3215
rect 1991 3231 1995 3235
rect 2024 3227 2028 3231
rect 1622 3171 1626 3175
rect 1632 3171 1636 3175
rect 1672 3173 1676 3177
rect 2109 3174 2113 3178
rect 2119 3174 2123 3178
rect 2159 3176 2163 3180
rect 1040 3130 1044 3134
rect 1050 3130 1054 3134
rect 1090 3132 1094 3136
rect 1155 3140 1159 3144
rect 1165 3140 1169 3144
rect 1205 3142 1209 3146
rect 1489 3118 1493 3122
rect 580 3086 584 3090
rect 596 3086 600 3090
rect 629 3082 633 3086
rect 684 3082 688 3086
rect 694 3082 698 3086
rect 734 3084 738 3088
rect 919 3095 923 3099
rect 1505 3118 1509 3122
rect 1538 3114 1542 3118
rect 935 3095 939 3099
rect 968 3091 972 3095
rect 1974 3103 1978 3107
rect 1990 3103 1994 3107
rect 2023 3099 2027 3103
rect 584 2982 588 2986
rect 629 2993 633 2997
rect 645 2993 649 2997
rect 678 2989 682 2993
rect 936 2984 940 2988
rect 981 2995 985 2999
rect 997 2995 1001 2999
rect 1030 2991 1034 2995
rect 1497 2984 1501 2989
rect 1542 2995 1546 2999
rect 2172 3003 2176 3007
rect 1558 2995 1562 2999
rect 1591 2991 1595 2995
rect 2217 3014 2221 3018
rect 2233 3014 2237 3018
rect 2266 3010 2270 3014
rect 737 2947 741 2951
rect 584 2926 588 2930
rect 631 2927 635 2931
rect 747 2947 751 2951
rect 787 2949 791 2953
rect 1089 2949 1093 2953
rect 647 2927 651 2931
rect 680 2923 684 2927
rect 936 2928 940 2932
rect 983 2929 987 2933
rect 1099 2949 1103 2953
rect 1139 2951 1143 2955
rect 1650 2949 1654 2953
rect 999 2929 1003 2933
rect 1032 2925 1036 2929
rect 1497 2928 1501 2932
rect 1544 2929 1548 2933
rect 1660 2949 1664 2953
rect 1700 2951 1704 2955
rect 2325 2968 2329 2972
rect 2172 2947 2176 2951
rect 2219 2948 2223 2952
rect 1560 2929 1564 2933
rect 1593 2925 1597 2929
rect 2335 2968 2339 2972
rect 2375 2970 2379 2974
rect 2235 2948 2239 2952
rect 2268 2944 2272 2948
rect 2206 2869 2210 2873
rect 2222 2869 2226 2873
rect 2255 2865 2259 2869
rect 986 2837 990 2842
rect 599 2817 603 2822
rect 1002 2838 1006 2842
rect 1035 2834 1039 2838
rect 1536 2838 1540 2843
rect 1552 2839 1556 2843
rect 1585 2835 1589 2839
rect 615 2818 619 2822
rect 648 2814 652 2818
<< metal1 >>
rect 2512 3899 2546 3903
rect 2518 3894 2522 3899
rect 2536 3894 2540 3899
rect 2560 3897 2594 3901
rect 2466 3890 2500 3894
rect 1890 3881 1924 3885
rect 2472 3884 2476 3890
rect 2566 3891 2570 3897
rect 1896 3876 1900 3881
rect 1914 3876 1918 3881
rect 1938 3879 1972 3883
rect 1844 3872 1878 3876
rect 1850 3866 1854 3872
rect 1944 3873 1948 3879
rect 1169 3855 1203 3859
rect 1759 3857 1829 3864
rect 1175 3850 1179 3855
rect 1193 3850 1197 3855
rect 1217 3853 1251 3857
rect 1123 3846 1157 3850
rect 1129 3840 1133 3846
rect 1223 3847 1227 3853
rect 1073 3833 1108 3838
rect 1073 3810 1078 3833
rect 1099 3822 1102 3823
rect 1147 3822 1151 3830
rect 1160 3829 1176 3833
rect 1160 3822 1164 3829
rect 1184 3826 1188 3840
rect 1196 3829 1200 3833
rect 1241 3829 1245 3837
rect 1184 3825 1197 3826
rect 1210 3825 1225 3829
rect 1241 3825 1261 3829
rect 1184 3822 1214 3825
rect 1241 3822 1245 3825
rect 1099 3818 1131 3822
rect 1147 3818 1164 3822
rect 1193 3821 1214 3822
rect 1147 3815 1151 3818
rect 391 3805 1078 3810
rect 1223 3811 1227 3817
rect 391 3345 396 3805
rect 1129 3804 1133 3810
rect 1175 3807 1179 3811
rect 1217 3808 1251 3811
rect 1169 3804 1203 3807
rect 1123 3801 1157 3804
rect 1123 3790 1157 3794
rect 1129 3784 1133 3790
rect 1171 3789 1205 3793
rect 1177 3784 1181 3789
rect 1195 3784 1199 3789
rect 1219 3787 1253 3791
rect 1256 3787 1261 3825
rect 1277 3822 1311 3826
rect 1283 3814 1287 3822
rect 1326 3813 1360 3817
rect 1332 3807 1336 3813
rect 1225 3781 1229 3787
rect 1256 3783 1284 3787
rect 1301 3781 1305 3794
rect 1350 3790 1354 3797
rect 1314 3785 1334 3789
rect 1350 3785 1367 3790
rect 1314 3781 1318 3785
rect 1350 3782 1354 3785
rect 1147 3766 1151 3774
rect 1161 3766 1178 3767
rect 1115 3762 1131 3766
rect 1147 3763 1178 3766
rect 1147 3762 1162 3763
rect 1147 3759 1151 3762
rect 1186 3760 1190 3774
rect 1301 3780 1318 3781
rect 1291 3777 1318 3780
rect 1291 3774 1297 3777
rect 1198 3763 1202 3767
rect 1243 3763 1247 3771
rect 1332 3771 1336 3777
rect 1186 3759 1199 3760
rect 1212 3759 1227 3763
rect 1243 3759 1257 3763
rect 1283 3763 1287 3769
rect 1301 3763 1305 3769
rect 1326 3768 1360 3771
rect 1277 3760 1311 3763
rect 1186 3756 1216 3759
rect 1243 3756 1247 3759
rect 1195 3755 1216 3756
rect 1129 3748 1133 3754
rect 1123 3745 1157 3748
rect 1225 3745 1229 3751
rect 1177 3741 1181 3745
rect 1219 3742 1253 3745
rect 1171 3738 1202 3741
rect 1759 3634 1768 3857
rect 1820 3848 1823 3849
rect 1868 3848 1872 3856
rect 1881 3855 1897 3859
rect 1881 3848 1885 3855
rect 1905 3852 1909 3866
rect 1917 3855 1921 3859
rect 1962 3855 1966 3863
rect 2442 3866 2445 3867
rect 2490 3866 2494 3874
rect 2503 3873 2519 3877
rect 2503 3866 2507 3873
rect 2527 3870 2531 3884
rect 2539 3873 2543 3877
rect 2584 3873 2588 3881
rect 2527 3869 2540 3870
rect 2553 3869 2568 3873
rect 2584 3869 2604 3873
rect 2527 3866 2557 3869
rect 2584 3866 2588 3869
rect 2442 3862 2474 3866
rect 2490 3862 2507 3866
rect 2536 3865 2557 3866
rect 2490 3859 2494 3862
rect 1905 3851 1918 3852
rect 1931 3851 1946 3855
rect 1962 3851 1982 3855
rect 2566 3855 2570 3861
rect 1905 3848 1935 3851
rect 1962 3848 1966 3851
rect 1820 3844 1852 3848
rect 1868 3844 1885 3848
rect 1914 3847 1935 3848
rect 1868 3841 1872 3844
rect 1944 3837 1948 3843
rect 1850 3830 1854 3836
rect 1896 3833 1900 3837
rect 1938 3834 1972 3837
rect 1890 3830 1924 3833
rect 1844 3827 1878 3830
rect 1844 3816 1878 3820
rect 1850 3810 1854 3816
rect 1892 3815 1926 3819
rect 1898 3810 1902 3815
rect 1916 3810 1920 3815
rect 1940 3813 1974 3817
rect 1977 3813 1982 3851
rect 1998 3848 2032 3852
rect 2472 3848 2476 3854
rect 2518 3851 2522 3855
rect 2560 3852 2594 3855
rect 2512 3848 2546 3851
rect 2004 3840 2008 3848
rect 2466 3845 2500 3848
rect 2047 3839 2081 3843
rect 2053 3833 2057 3839
rect 2466 3834 2500 3838
rect 1946 3807 1950 3813
rect 1977 3809 2005 3813
rect 2022 3807 2026 3820
rect 2071 3816 2075 3823
rect 2472 3828 2476 3834
rect 2514 3833 2548 3837
rect 2520 3828 2524 3833
rect 2538 3828 2542 3833
rect 2562 3831 2596 3835
rect 2599 3831 2604 3869
rect 2620 3866 2654 3870
rect 2626 3858 2630 3866
rect 2669 3857 2703 3861
rect 2675 3851 2679 3857
rect 2568 3825 2572 3831
rect 2599 3827 2627 3831
rect 2644 3825 2648 3838
rect 2693 3834 2697 3841
rect 2657 3829 2677 3833
rect 2693 3829 2716 3834
rect 2657 3825 2661 3829
rect 2693 3826 2697 3829
rect 2035 3811 2055 3815
rect 2071 3811 2092 3816
rect 2035 3807 2039 3811
rect 2071 3808 2075 3811
rect 1868 3792 1872 3800
rect 1882 3792 1899 3793
rect 1836 3788 1852 3792
rect 1868 3789 1899 3792
rect 1868 3788 1883 3789
rect 1868 3785 1872 3788
rect 1907 3786 1911 3800
rect 2022 3806 2039 3807
rect 2012 3803 2039 3806
rect 2490 3810 2494 3818
rect 2504 3810 2521 3811
rect 2458 3806 2474 3810
rect 2490 3807 2521 3810
rect 2490 3806 2505 3807
rect 2490 3803 2494 3806
rect 2012 3800 2018 3803
rect 1919 3789 1923 3793
rect 1964 3789 1968 3797
rect 2053 3797 2057 3803
rect 2529 3804 2533 3818
rect 2644 3824 2661 3825
rect 2634 3821 2661 3824
rect 2634 3818 2640 3821
rect 2675 3815 2679 3821
rect 2541 3807 2545 3811
rect 2626 3807 2630 3813
rect 2644 3807 2648 3813
rect 2669 3812 2703 3815
rect 2529 3803 2542 3804
rect 2555 3803 2570 3807
rect 2620 3804 2654 3807
rect 2529 3800 2559 3803
rect 2538 3799 2559 3800
rect 1907 3785 1920 3786
rect 1933 3785 1948 3789
rect 1964 3785 1978 3789
rect 2004 3789 2008 3795
rect 2022 3789 2026 3795
rect 2047 3794 2081 3797
rect 2472 3792 2476 3798
rect 2466 3789 2500 3792
rect 2568 3789 2572 3795
rect 1998 3786 2032 3789
rect 2520 3785 2524 3789
rect 2562 3786 2596 3789
rect 1907 3782 1937 3785
rect 1964 3782 1968 3785
rect 2514 3782 2545 3785
rect 1916 3781 1937 3782
rect 1850 3774 1854 3780
rect 1844 3771 1878 3774
rect 1946 3771 1950 3777
rect 1898 3767 1902 3771
rect 1940 3768 1974 3771
rect 1892 3764 1923 3767
rect 1391 3630 1768 3634
rect 1248 3629 1767 3630
rect 1248 3625 1396 3629
rect 624 3609 658 3613
rect 630 3604 634 3609
rect 648 3604 652 3609
rect 672 3607 706 3611
rect 578 3600 612 3604
rect 584 3594 588 3600
rect 678 3601 682 3607
rect 467 3345 472 3584
rect 554 3576 557 3577
rect 602 3576 606 3584
rect 615 3583 631 3587
rect 615 3576 619 3583
rect 639 3580 643 3594
rect 651 3583 655 3587
rect 696 3583 700 3591
rect 639 3579 652 3580
rect 665 3579 680 3583
rect 696 3579 716 3583
rect 639 3576 669 3579
rect 696 3576 700 3579
rect 554 3572 586 3576
rect 602 3572 619 3576
rect 648 3575 669 3576
rect 602 3569 606 3572
rect 678 3565 682 3571
rect 584 3558 588 3564
rect 630 3561 634 3565
rect 672 3562 706 3565
rect 624 3558 658 3561
rect 578 3555 612 3558
rect 578 3544 612 3548
rect 584 3538 588 3544
rect 626 3543 660 3547
rect 632 3538 636 3543
rect 650 3538 654 3543
rect 674 3541 708 3545
rect 711 3541 716 3579
rect 732 3576 766 3580
rect 738 3568 742 3576
rect 781 3567 815 3571
rect 787 3561 791 3567
rect 680 3535 684 3541
rect 711 3537 739 3541
rect 756 3535 760 3548
rect 805 3544 809 3551
rect 769 3539 789 3543
rect 805 3539 851 3544
rect 769 3535 773 3539
rect 805 3536 809 3539
rect 602 3520 606 3528
rect 616 3520 633 3521
rect 570 3516 586 3520
rect 602 3517 633 3520
rect 602 3516 617 3517
rect 602 3513 606 3516
rect 641 3514 645 3528
rect 756 3534 773 3535
rect 746 3531 773 3534
rect 746 3528 752 3531
rect 653 3517 657 3521
rect 698 3517 702 3525
rect 787 3525 791 3531
rect 641 3513 654 3514
rect 667 3513 682 3517
rect 698 3513 712 3517
rect 738 3517 742 3523
rect 756 3517 760 3523
rect 781 3522 815 3525
rect 732 3514 766 3517
rect 641 3510 671 3513
rect 698 3510 702 3513
rect 650 3509 671 3510
rect 584 3502 588 3508
rect 578 3499 612 3502
rect 680 3499 684 3505
rect 632 3495 636 3499
rect 674 3496 708 3499
rect 626 3492 657 3495
rect 391 2706 396 3338
rect 467 2780 472 3338
rect 907 3230 941 3234
rect 913 3225 917 3230
rect 931 3225 935 3230
rect 955 3228 989 3232
rect 961 3222 965 3228
rect 899 3203 914 3208
rect 922 3201 926 3215
rect 922 3200 935 3201
rect 944 3200 963 3204
rect 922 3197 947 3200
rect 931 3196 947 3197
rect 961 3186 965 3192
rect 913 3182 917 3186
rect 955 3183 989 3186
rect 907 3179 941 3182
rect 1148 3179 1182 3183
rect 1033 3169 1067 3173
rect 1154 3171 1158 3179
rect 1039 3161 1043 3169
rect 1082 3160 1116 3164
rect 1088 3154 1092 3160
rect 1197 3170 1231 3174
rect 1203 3164 1207 3170
rect 665 3128 905 3132
rect 573 3112 607 3116
rect 579 3107 583 3112
rect 597 3107 601 3112
rect 621 3110 655 3114
rect 627 3104 631 3110
rect 554 3086 580 3090
rect 554 3039 560 3086
rect 588 3083 592 3097
rect 645 3086 649 3094
rect 665 3086 669 3128
rect 677 3121 711 3125
rect 683 3113 687 3121
rect 726 3112 760 3116
rect 732 3106 736 3112
rect 588 3082 601 3083
rect 610 3082 629 3086
rect 645 3082 684 3086
rect 588 3079 613 3082
rect 645 3079 649 3082
rect 701 3080 705 3093
rect 750 3089 754 3096
rect 900 3099 905 3128
rect 1057 3128 1061 3141
rect 1106 3136 1110 3144
rect 1117 3140 1155 3144
rect 1117 3136 1121 3140
rect 1172 3138 1176 3151
rect 1221 3146 1225 3154
rect 1248 3146 1253 3625
rect 1571 3507 1942 3512
rect 1479 3347 1513 3351
rect 1485 3342 1489 3347
rect 1503 3342 1507 3347
rect 1527 3345 1561 3349
rect 1533 3339 1537 3345
rect 1450 3321 1486 3325
rect 1450 3219 1456 3321
rect 1494 3318 1498 3332
rect 1551 3321 1555 3329
rect 1571 3321 1577 3507
rect 1964 3503 1998 3507
rect 1970 3498 1974 3503
rect 1988 3498 1992 3503
rect 2012 3501 2046 3505
rect 2018 3495 2022 3501
rect 1920 3476 1932 3481
rect 1937 3476 1971 3481
rect 1920 3358 1924 3476
rect 1979 3474 1983 3488
rect 2036 3477 2040 3485
rect 1979 3473 1992 3474
rect 2001 3473 2020 3477
rect 2036 3473 2059 3477
rect 1979 3470 2004 3473
rect 2036 3470 2040 3473
rect 1988 3469 2004 3470
rect 2018 3459 2022 3465
rect 1970 3455 1974 3459
rect 2012 3456 2046 3459
rect 1964 3452 1998 3455
rect 2056 3422 2059 3473
rect 2103 3457 2137 3461
rect 2109 3449 2113 3457
rect 2152 3448 2186 3452
rect 2158 3442 2162 3448
rect 2056 3418 2110 3422
rect 2127 3416 2131 3429
rect 2176 3424 2180 3432
rect 2140 3420 2160 3424
rect 2176 3420 2240 3424
rect 2140 3416 2144 3420
rect 2176 3417 2180 3420
rect 2127 3415 2144 3416
rect 2117 3412 2144 3415
rect 2117 3409 2123 3412
rect 2158 3406 2162 3412
rect 2109 3398 2113 3404
rect 2127 3398 2131 3404
rect 2152 3403 2186 3406
rect 2103 3395 2137 3398
rect 1963 3380 1997 3384
rect 1969 3375 1973 3380
rect 1987 3375 1991 3380
rect 2011 3378 2045 3382
rect 2017 3372 2021 3378
rect 1920 3354 1970 3358
rect 1494 3317 1507 3318
rect 1516 3317 1535 3321
rect 1551 3317 1587 3321
rect 1494 3314 1519 3317
rect 1551 3314 1555 3317
rect 1503 3313 1519 3314
rect 1533 3303 1537 3309
rect 1485 3299 1489 3303
rect 1527 3300 1561 3303
rect 1479 3296 1513 3299
rect 1583 3277 1587 3317
rect 1611 3312 1645 3316
rect 1617 3304 1621 3312
rect 1660 3303 1694 3307
rect 1666 3297 1670 3303
rect 1583 3273 1618 3277
rect 1635 3271 1639 3284
rect 1684 3279 1688 3287
rect 1648 3275 1668 3279
rect 1684 3275 1704 3279
rect 1648 3271 1652 3275
rect 1684 3272 1688 3275
rect 1635 3270 1652 3271
rect 1625 3267 1652 3270
rect 1625 3264 1631 3267
rect 1666 3261 1670 3267
rect 1617 3253 1621 3259
rect 1635 3253 1639 3259
rect 1660 3258 1694 3261
rect 1611 3250 1645 3253
rect 1478 3241 1512 3245
rect 1484 3236 1488 3241
rect 1502 3236 1506 3241
rect 1526 3239 1560 3243
rect 1532 3233 1536 3239
rect 1701 3238 1704 3275
rect 1727 3273 1761 3277
rect 1733 3265 1737 3273
rect 1776 3264 1810 3268
rect 1782 3258 1786 3264
rect 1701 3234 1734 3238
rect 1450 3215 1485 3219
rect 1450 3175 1456 3215
rect 1493 3212 1497 3226
rect 1751 3232 1755 3245
rect 1800 3240 1804 3248
rect 1764 3236 1784 3240
rect 1800 3236 1812 3240
rect 1764 3232 1768 3236
rect 1800 3233 1804 3236
rect 1751 3231 1768 3232
rect 1741 3228 1768 3231
rect 1741 3225 1747 3228
rect 1782 3222 1786 3228
rect 1493 3211 1506 3212
rect 1515 3211 1534 3215
rect 1733 3214 1737 3220
rect 1751 3214 1755 3220
rect 1776 3219 1810 3222
rect 1493 3208 1518 3211
rect 1615 3210 1649 3214
rect 1727 3211 1761 3214
rect 1502 3207 1518 3208
rect 1532 3197 1536 3203
rect 1621 3202 1625 3210
rect 1484 3193 1488 3197
rect 1526 3194 1560 3197
rect 1478 3190 1512 3193
rect 1664 3201 1698 3205
rect 1670 3195 1674 3201
rect 1450 3169 1587 3175
rect 1185 3142 1205 3146
rect 1221 3142 1253 3146
rect 1482 3144 1516 3148
rect 1185 3138 1189 3142
rect 1221 3139 1225 3142
rect 1172 3137 1189 3138
rect 1070 3132 1090 3136
rect 1106 3132 1121 3136
rect 1162 3134 1189 3137
rect 1488 3139 1492 3144
rect 1506 3139 1510 3144
rect 1530 3142 1564 3146
rect 1070 3128 1074 3132
rect 1106 3129 1110 3132
rect 1162 3131 1168 3134
rect 1057 3127 1074 3128
rect 912 3121 946 3125
rect 1047 3124 1074 3127
rect 1203 3128 1207 3134
rect 1536 3136 1540 3142
rect 918 3116 922 3121
rect 936 3116 940 3121
rect 960 3119 994 3123
rect 1047 3121 1053 3124
rect 966 3113 970 3119
rect 1088 3118 1092 3124
rect 1154 3120 1158 3126
rect 1172 3120 1176 3126
rect 1197 3125 1231 3128
rect 900 3095 919 3099
rect 927 3092 931 3106
rect 1039 3110 1043 3116
rect 1057 3110 1061 3116
rect 1082 3115 1116 3118
rect 1148 3117 1182 3120
rect 1459 3118 1489 3122
rect 1033 3107 1067 3110
rect 984 3095 988 3103
rect 927 3091 940 3092
rect 949 3091 968 3095
rect 984 3091 1021 3095
rect 714 3084 734 3088
rect 750 3084 769 3089
rect 927 3088 952 3091
rect 984 3088 988 3091
rect 936 3087 952 3088
rect 714 3080 718 3084
rect 750 3081 754 3084
rect 701 3079 718 3080
rect 597 3078 613 3079
rect 691 3076 718 3079
rect 966 3077 970 3083
rect 627 3068 631 3074
rect 691 3073 697 3076
rect 732 3070 736 3076
rect 918 3073 922 3077
rect 960 3074 994 3077
rect 912 3070 946 3073
rect 579 3064 583 3068
rect 621 3065 655 3068
rect 573 3061 607 3064
rect 683 3062 687 3068
rect 701 3062 705 3068
rect 726 3067 760 3070
rect 677 3059 711 3062
rect 862 3054 1145 3062
rect 554 3032 822 3039
rect 622 3019 656 3023
rect 628 3014 632 3019
rect 646 3014 650 3019
rect 670 3017 704 3021
rect 576 3010 610 3014
rect 582 3004 586 3010
rect 676 3011 680 3017
rect 552 2986 555 2987
rect 600 2986 604 2994
rect 613 2993 629 2997
rect 613 2986 617 2993
rect 637 2990 641 3004
rect 649 2993 653 2997
rect 694 2993 698 3001
rect 637 2989 650 2990
rect 663 2989 678 2993
rect 694 2989 714 2993
rect 637 2986 667 2989
rect 694 2986 698 2989
rect 552 2982 584 2986
rect 600 2982 617 2986
rect 646 2985 667 2986
rect 600 2979 604 2982
rect 676 2975 680 2981
rect 582 2968 586 2974
rect 628 2971 632 2975
rect 670 2972 704 2975
rect 622 2968 656 2971
rect 576 2965 610 2968
rect 576 2954 610 2958
rect 582 2948 586 2954
rect 624 2953 658 2957
rect 630 2948 634 2953
rect 648 2948 652 2953
rect 672 2951 706 2955
rect 709 2951 714 2989
rect 730 2986 764 2990
rect 736 2978 740 2986
rect 779 2977 813 2981
rect 785 2971 789 2977
rect 678 2945 682 2951
rect 709 2947 737 2951
rect 754 2945 758 2958
rect 803 2953 807 2961
rect 818 2953 822 3032
rect 767 2949 787 2953
rect 803 2949 822 2953
rect 767 2945 771 2949
rect 803 2946 807 2949
rect 600 2930 604 2938
rect 614 2930 631 2931
rect 568 2926 584 2930
rect 600 2927 631 2930
rect 600 2926 615 2927
rect 600 2923 604 2926
rect 639 2924 643 2938
rect 754 2944 771 2945
rect 744 2941 771 2944
rect 744 2938 750 2941
rect 651 2927 655 2931
rect 696 2927 700 2935
rect 785 2935 789 2941
rect 639 2923 652 2924
rect 665 2923 680 2927
rect 696 2923 710 2927
rect 736 2927 740 2933
rect 754 2927 758 2933
rect 779 2932 813 2935
rect 730 2924 764 2927
rect 639 2920 669 2923
rect 696 2920 700 2923
rect 648 2919 669 2920
rect 582 2912 586 2918
rect 576 2909 610 2912
rect 678 2909 682 2915
rect 630 2905 634 2909
rect 672 2906 706 2909
rect 624 2902 655 2905
rect 592 2844 626 2848
rect 598 2839 602 2844
rect 616 2839 620 2844
rect 640 2842 674 2846
rect 646 2836 650 2842
rect 590 2817 599 2822
rect 607 2815 611 2829
rect 664 2818 668 2826
rect 607 2814 620 2815
rect 629 2814 648 2818
rect 607 2811 632 2814
rect 664 2813 678 2818
rect 664 2811 668 2813
rect 616 2810 632 2811
rect 646 2800 650 2806
rect 598 2796 602 2800
rect 640 2797 674 2800
rect 592 2793 626 2796
rect 818 2780 822 2949
rect 863 2807 868 3054
rect 974 3021 1008 3025
rect 980 3016 984 3021
rect 998 3016 1002 3021
rect 1022 3019 1056 3023
rect 928 3012 962 3016
rect 934 3006 938 3012
rect 1028 3013 1032 3019
rect 904 2988 907 2989
rect 952 2988 956 2996
rect 965 2995 981 2999
rect 965 2988 969 2995
rect 989 2992 993 3006
rect 1001 2995 1005 2999
rect 1046 2995 1050 3003
rect 989 2991 1002 2992
rect 1015 2991 1030 2995
rect 1046 2991 1066 2995
rect 989 2988 1019 2991
rect 1046 2988 1050 2991
rect 904 2984 936 2988
rect 952 2984 969 2988
rect 998 2987 1019 2988
rect 952 2981 956 2984
rect 1028 2977 1032 2983
rect 934 2970 938 2976
rect 980 2973 984 2977
rect 1022 2974 1056 2977
rect 974 2970 1008 2973
rect 928 2967 962 2970
rect 928 2956 962 2960
rect 934 2950 938 2956
rect 976 2955 1010 2959
rect 982 2950 986 2955
rect 1000 2950 1004 2955
rect 1024 2953 1058 2957
rect 1061 2953 1066 2991
rect 1082 2988 1116 2992
rect 1088 2980 1092 2988
rect 1170 2983 1175 3051
rect 1131 2979 1165 2983
rect 1137 2973 1141 2979
rect 1030 2947 1034 2953
rect 1061 2949 1089 2953
rect 1106 2947 1110 2960
rect 1155 2955 1159 2963
rect 1170 2955 1175 2978
rect 1119 2951 1139 2955
rect 1155 2951 1175 2955
rect 1119 2947 1123 2951
rect 1155 2948 1159 2951
rect 952 2932 956 2940
rect 966 2932 983 2933
rect 920 2928 936 2932
rect 952 2929 983 2932
rect 952 2928 967 2929
rect 952 2925 956 2928
rect 991 2926 995 2940
rect 1106 2946 1123 2947
rect 1096 2943 1123 2946
rect 1096 2940 1102 2943
rect 1003 2929 1007 2933
rect 1048 2929 1052 2937
rect 1137 2937 1141 2943
rect 991 2925 1004 2926
rect 1017 2925 1032 2929
rect 1048 2925 1062 2929
rect 1088 2929 1092 2935
rect 1106 2929 1110 2935
rect 1131 2934 1165 2937
rect 1082 2926 1116 2929
rect 991 2922 1021 2925
rect 1048 2922 1052 2925
rect 1000 2921 1021 2922
rect 934 2914 938 2920
rect 928 2911 962 2914
rect 1030 2911 1034 2917
rect 982 2907 986 2911
rect 1024 2908 1058 2911
rect 976 2904 1007 2907
rect 979 2864 1013 2868
rect 985 2859 989 2864
rect 1003 2859 1007 2864
rect 1027 2862 1061 2866
rect 1033 2856 1037 2862
rect 944 2837 986 2842
rect 994 2835 998 2849
rect 1051 2838 1055 2846
rect 994 2834 1007 2835
rect 1016 2834 1035 2838
rect 1051 2834 1086 2838
rect 994 2831 1019 2834
rect 1051 2831 1055 2834
rect 1003 2830 1019 2831
rect 1082 2829 1086 2834
rect 1220 2829 1225 3072
rect 1459 3053 1465 3118
rect 1497 3115 1501 3129
rect 1497 3114 1510 3115
rect 1519 3114 1538 3118
rect 1497 3111 1522 3114
rect 1506 3110 1522 3111
rect 1536 3100 1540 3106
rect 1488 3096 1492 3100
rect 1530 3097 1564 3100
rect 1482 3093 1516 3096
rect 1579 3053 1587 3169
rect 1599 3171 1622 3175
rect 1599 3074 1605 3171
rect 1639 3169 1643 3182
rect 1652 3173 1672 3177
rect 1652 3169 1656 3173
rect 1639 3168 1656 3169
rect 1629 3165 1656 3168
rect 1629 3162 1635 3165
rect 1670 3159 1674 3165
rect 1621 3151 1625 3157
rect 1639 3151 1643 3157
rect 1664 3156 1698 3159
rect 1615 3148 1649 3151
rect 1845 3074 1850 3261
rect 1599 3065 1850 3074
rect 1920 3235 1924 3354
rect 1978 3351 1982 3365
rect 1978 3350 1991 3351
rect 2000 3350 2019 3354
rect 1978 3347 2003 3350
rect 1987 3346 2003 3347
rect 2017 3336 2021 3342
rect 1969 3332 1973 3336
rect 2011 3333 2045 3336
rect 1963 3329 1997 3332
rect 2236 3302 2240 3420
rect 2464 3346 2498 3350
rect 2279 3337 2313 3341
rect 2470 3338 2474 3346
rect 2285 3329 2289 3337
rect 2328 3328 2362 3332
rect 2334 3322 2338 3328
rect 2513 3337 2547 3341
rect 2519 3331 2523 3337
rect 2236 3298 2286 3302
rect 2303 3296 2307 3309
rect 2352 3304 2356 3312
rect 2398 3307 2471 3311
rect 2398 3304 2402 3307
rect 2488 3305 2492 3318
rect 2501 3309 2521 3313
rect 2501 3305 2505 3309
rect 2488 3304 2505 3305
rect 2316 3300 2336 3304
rect 2352 3300 2402 3304
rect 2478 3301 2505 3304
rect 2316 3296 2320 3300
rect 2352 3297 2356 3300
rect 2478 3298 2484 3301
rect 2303 3295 2320 3296
rect 2293 3292 2320 3295
rect 2519 3295 2523 3301
rect 2293 3289 2299 3292
rect 2334 3286 2338 3292
rect 2470 3287 2474 3293
rect 2488 3287 2492 3293
rect 2513 3292 2547 3295
rect 2285 3278 2289 3284
rect 2303 3278 2307 3284
rect 2328 3283 2362 3286
rect 2464 3284 2498 3287
rect 2279 3275 2313 3278
rect 1968 3257 2002 3261
rect 1974 3252 1978 3257
rect 1992 3252 1996 3257
rect 2016 3255 2050 3259
rect 2022 3249 2026 3255
rect 1920 3231 1975 3235
rect 1920 3107 1924 3231
rect 1983 3228 1987 3242
rect 2040 3231 2044 3239
rect 1983 3227 1996 3228
rect 2005 3227 2024 3231
rect 2040 3227 2063 3231
rect 1983 3224 2008 3227
rect 2040 3224 2044 3227
rect 1992 3223 2008 3224
rect 2022 3213 2026 3219
rect 1974 3209 1978 3213
rect 2016 3210 2050 3213
rect 1968 3206 2002 3209
rect 2060 3178 2063 3227
rect 2102 3213 2136 3217
rect 2108 3205 2112 3213
rect 2151 3204 2185 3208
rect 2157 3198 2161 3204
rect 2060 3174 2109 3178
rect 2126 3172 2130 3185
rect 2139 3176 2159 3180
rect 2139 3172 2143 3176
rect 2126 3171 2143 3172
rect 2116 3168 2143 3171
rect 2116 3165 2122 3168
rect 2157 3162 2161 3168
rect 2108 3154 2112 3160
rect 2126 3154 2130 3160
rect 2151 3159 2185 3162
rect 2102 3151 2136 3154
rect 1967 3129 2001 3133
rect 1973 3124 1977 3129
rect 1991 3124 1995 3129
rect 2015 3127 2049 3131
rect 2021 3121 2025 3127
rect 1920 3103 1974 3107
rect 1920 3072 1924 3103
rect 1982 3100 1986 3114
rect 1982 3099 1995 3100
rect 2004 3099 2023 3103
rect 1982 3096 2007 3099
rect 1991 3095 2007 3096
rect 2021 3085 2025 3091
rect 1973 3081 1977 3085
rect 2015 3082 2049 3085
rect 1967 3078 2001 3081
rect 1920 3066 2410 3072
rect 1459 3048 1735 3053
rect 1535 3021 1569 3025
rect 1541 3016 1545 3021
rect 1559 3016 1563 3021
rect 1583 3019 1617 3023
rect 1489 3012 1523 3016
rect 1495 3006 1499 3012
rect 1589 3013 1593 3019
rect 1465 2984 1497 2989
rect 1513 2988 1517 2996
rect 1526 2995 1542 2999
rect 1526 2988 1530 2995
rect 1550 2992 1554 3006
rect 1562 2995 1566 2999
rect 1607 2995 1611 3003
rect 1550 2991 1563 2992
rect 1576 2991 1591 2995
rect 1607 2991 1627 2995
rect 1550 2988 1580 2991
rect 1607 2988 1611 2991
rect 1513 2984 1530 2988
rect 1559 2987 1580 2988
rect 1033 2820 1037 2826
rect 1082 2825 1225 2829
rect 1513 2981 1517 2984
rect 985 2816 989 2820
rect 1027 2817 1061 2820
rect 979 2813 1013 2816
rect 1082 2807 1086 2825
rect 863 2802 1086 2807
rect 467 2776 822 2780
rect 1264 2706 1269 2978
rect 1589 2977 1593 2983
rect 1495 2970 1499 2976
rect 1541 2973 1545 2977
rect 1583 2974 1617 2977
rect 1535 2970 1569 2973
rect 1489 2967 1523 2970
rect 1489 2956 1523 2960
rect 1495 2950 1499 2956
rect 1537 2955 1571 2959
rect 1543 2950 1547 2955
rect 1561 2950 1565 2955
rect 1585 2953 1619 2957
rect 1622 2953 1627 2991
rect 1643 2988 1677 2992
rect 1649 2980 1653 2988
rect 1692 2979 1726 2983
rect 1698 2973 1702 2979
rect 1591 2947 1595 2953
rect 1622 2949 1650 2953
rect 1667 2947 1671 2960
rect 1716 2955 1720 2963
rect 1730 2956 1735 3048
rect 1680 2951 1700 2955
rect 1716 2951 1730 2955
rect 1680 2947 1684 2951
rect 1716 2948 1720 2951
rect 1513 2932 1517 2940
rect 1527 2932 1544 2933
rect 1481 2928 1497 2932
rect 1513 2929 1544 2932
rect 1513 2928 1528 2929
rect 1513 2925 1517 2928
rect 1552 2926 1556 2940
rect 1667 2946 1684 2947
rect 1657 2943 1684 2946
rect 1657 2940 1663 2943
rect 1564 2929 1568 2933
rect 1609 2929 1613 2937
rect 1698 2937 1702 2943
rect 1552 2925 1565 2926
rect 1578 2925 1593 2929
rect 1609 2925 1623 2929
rect 1649 2929 1653 2935
rect 1667 2929 1671 2935
rect 1692 2934 1726 2937
rect 1643 2926 1677 2929
rect 1552 2922 1582 2925
rect 1609 2922 1613 2925
rect 1561 2921 1582 2922
rect 1495 2914 1499 2920
rect 1489 2911 1523 2914
rect 1591 2911 1595 2917
rect 1543 2907 1547 2911
rect 1585 2908 1619 2911
rect 1537 2904 1568 2907
rect 1529 2865 1563 2869
rect 1535 2860 1539 2865
rect 1553 2860 1557 2865
rect 1577 2863 1611 2867
rect 1583 2857 1587 2863
rect 1505 2838 1536 2843
rect 1544 2836 1548 2850
rect 1601 2839 1605 2847
rect 1795 2839 1803 3065
rect 2210 3040 2244 3044
rect 2216 3035 2220 3040
rect 2234 3035 2238 3040
rect 2258 3038 2292 3042
rect 2164 3031 2198 3035
rect 2170 3025 2174 3031
rect 2264 3032 2268 3038
rect 2140 3007 2143 3008
rect 2188 3007 2192 3015
rect 2201 3014 2217 3018
rect 2201 3007 2205 3014
rect 2225 3011 2229 3025
rect 2237 3014 2241 3018
rect 2282 3014 2286 3022
rect 2225 3010 2238 3011
rect 2251 3010 2266 3014
rect 2282 3010 2302 3014
rect 2225 3007 2255 3010
rect 2282 3007 2286 3010
rect 2140 3003 2172 3007
rect 2188 3003 2205 3007
rect 2234 3006 2255 3007
rect 2188 3000 2192 3003
rect 2264 2996 2268 3002
rect 2170 2989 2174 2995
rect 2216 2992 2220 2996
rect 2258 2993 2292 2996
rect 2210 2989 2244 2992
rect 2164 2986 2198 2989
rect 2164 2975 2198 2979
rect 2170 2969 2174 2975
rect 2212 2974 2246 2978
rect 2218 2969 2222 2974
rect 2236 2969 2240 2974
rect 2260 2972 2294 2976
rect 2297 2972 2302 3010
rect 2318 3007 2352 3011
rect 2324 2999 2328 3007
rect 2367 2998 2401 3002
rect 2373 2992 2377 2998
rect 2266 2966 2270 2972
rect 2297 2968 2325 2972
rect 2342 2966 2346 2979
rect 2391 2974 2395 2982
rect 2406 2974 2410 3066
rect 2355 2970 2375 2974
rect 2391 2970 2410 2974
rect 2355 2966 2359 2970
rect 2391 2967 2395 2970
rect 2188 2951 2192 2959
rect 2202 2951 2219 2952
rect 2156 2947 2172 2951
rect 2188 2948 2219 2951
rect 2188 2947 2203 2948
rect 2149 2873 2156 2947
rect 2188 2944 2192 2947
rect 2227 2945 2231 2959
rect 2342 2965 2359 2966
rect 2332 2962 2359 2965
rect 2332 2959 2338 2962
rect 2373 2956 2377 2962
rect 2239 2948 2243 2952
rect 2324 2948 2328 2954
rect 2342 2948 2346 2954
rect 2367 2953 2401 2956
rect 2227 2944 2240 2945
rect 2253 2944 2268 2948
rect 2318 2945 2352 2948
rect 2227 2941 2257 2944
rect 2236 2940 2257 2941
rect 2170 2933 2174 2939
rect 2164 2930 2198 2933
rect 2266 2930 2270 2936
rect 2218 2926 2222 2930
rect 2260 2927 2294 2930
rect 2212 2923 2243 2926
rect 2199 2895 2233 2899
rect 2205 2890 2209 2895
rect 2223 2890 2227 2895
rect 2247 2893 2281 2897
rect 2253 2887 2257 2893
rect 2149 2869 2206 2873
rect 2214 2866 2218 2880
rect 2214 2865 2227 2866
rect 2236 2865 2255 2869
rect 2214 2862 2239 2865
rect 2223 2861 2239 2862
rect 2253 2851 2257 2857
rect 2205 2847 2209 2851
rect 2247 2848 2281 2851
rect 2199 2844 2233 2847
rect 1544 2835 1557 2836
rect 1566 2835 1585 2839
rect 1601 2835 1803 2839
rect 1544 2832 1569 2835
rect 1601 2832 1605 2835
rect 1553 2831 1569 2832
rect 1583 2821 1587 2827
rect 1535 2817 1539 2821
rect 1577 2818 1611 2821
rect 1529 2814 1563 2817
rect 391 2699 1269 2706
<< m2contact >>
rect 1829 3857 1836 3864
rect 1108 3833 1115 3838
rect 1094 3818 1099 3823
rect 1200 3828 1205 3833
rect 1367 3785 1374 3790
rect 1108 3762 1115 3767
rect 1202 3762 1207 3767
rect 1257 3759 1262 3764
rect 1815 3844 1820 3849
rect 1921 3854 1926 3859
rect 2437 3862 2442 3867
rect 2543 3872 2548 3877
rect 2716 3829 2722 3834
rect 2092 3811 2097 3816
rect 1829 3788 1836 3793
rect 2451 3806 2458 3811
rect 1923 3788 1928 3793
rect 2545 3806 2550 3811
rect 1978 3785 1983 3790
rect 467 3584 472 3589
rect 549 3572 554 3577
rect 655 3582 660 3587
rect 851 3539 860 3544
rect 563 3516 570 3521
rect 657 3516 662 3521
rect 712 3513 717 3518
rect 894 3203 899 3208
rect 1942 3507 1947 3512
rect 1932 3476 1937 3481
rect 1845 3261 1850 3266
rect 1812 3236 1817 3241
rect 1015 3095 1021 3100
rect 769 3084 774 3089
rect 1220 3072 1225 3077
rect 1137 3062 1145 3069
rect 547 2982 552 2987
rect 653 2992 658 2997
rect 561 2926 568 2931
rect 655 2926 660 2931
rect 710 2923 715 2928
rect 585 2817 590 2822
rect 678 2813 683 2818
rect 1163 3044 1170 3051
rect 899 2984 904 2989
rect 1005 2994 1010 2999
rect 1170 2978 1175 2983
rect 913 2928 920 2933
rect 1007 2928 1012 2933
rect 1062 2925 1067 2930
rect 939 2837 944 2842
rect 1458 2984 1465 2989
rect 1566 2994 1571 2999
rect 1264 2978 1269 2983
rect 1730 2951 1735 2956
rect 1474 2928 1481 2933
rect 1568 2928 1573 2933
rect 1623 2925 1628 2930
rect 1500 2838 1505 2843
rect 2135 3003 2140 3008
rect 2241 3013 2246 3018
rect 2149 2947 2156 2952
rect 2243 2947 2248 2952
<< metal2 >>
rect 563 3617 664 3621
rect 563 3589 570 3617
rect 472 3584 570 3589
rect 549 3491 554 3572
rect 563 3521 570 3584
rect 660 3582 664 3617
rect 851 3544 860 3930
rect 1108 3863 1209 3867
rect 1108 3838 1115 3863
rect 1094 3751 1099 3818
rect 1108 3767 1115 3833
rect 1205 3828 1209 3863
rect 1367 3790 1374 3930
rect 1829 3889 1930 3893
rect 1829 3864 1836 3889
rect 1292 3783 1298 3787
rect 1257 3780 1295 3783
rect 1094 3737 1099 3741
rect 1202 3737 1207 3762
rect 1257 3764 1262 3780
rect 1815 3763 1820 3844
rect 1829 3793 1836 3857
rect 1926 3854 1930 3889
rect 2092 3816 2097 3930
rect 2451 3907 2552 3911
rect 2451 3900 2458 3907
rect 2434 3862 2437 3867
rect 2434 3850 2442 3862
rect 2012 3809 2015 3813
rect 2377 3845 2442 3850
rect 1978 3806 2015 3809
rect 1923 3763 1928 3788
rect 1978 3790 1983 3806
rect 1815 3757 1867 3763
rect 1873 3757 1928 3763
rect 2377 3749 2381 3845
rect 2434 3781 2442 3845
rect 2451 3811 2458 3895
rect 2548 3872 2552 3907
rect 2716 3834 2722 3930
rect 2634 3827 2637 3831
rect 2600 3824 2637 3827
rect 2545 3781 2550 3806
rect 2586 3807 2590 3815
rect 2600 3807 2605 3824
rect 2586 3803 2605 3807
rect 2586 3800 2590 3803
rect 2434 3776 2550 3781
rect 1094 3731 1207 3737
rect 2056 3745 2381 3749
rect 746 3537 749 3541
rect 712 3534 749 3537
rect 657 3491 662 3516
rect 712 3518 717 3534
rect 2056 3529 2059 3745
rect 1932 3525 2059 3529
rect 555 3485 662 3491
rect 1932 3481 1937 3525
rect 1947 3507 2005 3512
rect 2001 3481 2005 3507
rect 1991 3477 2005 3481
rect 2117 3418 2120 3422
rect 2056 3415 2120 3418
rect 1592 3384 2004 3388
rect 1592 3273 1595 3384
rect 2000 3358 2004 3384
rect 1990 3354 2004 3358
rect 2035 3353 2039 3362
rect 2056 3353 2059 3415
rect 2035 3350 2059 3353
rect 2035 3347 2039 3350
rect 2537 3313 2541 3321
rect 2478 3307 2481 3311
rect 2425 3304 2481 3307
rect 2537 3309 2560 3313
rect 2537 3306 2541 3309
rect 2293 3298 2296 3302
rect 2264 3295 2296 3298
rect 1625 3273 1628 3277
rect 1569 3270 1628 3273
rect 945 3234 1008 3238
rect 945 3208 949 3234
rect 644 3203 894 3208
rect 934 3204 949 3208
rect 644 3132 649 3203
rect 1003 3133 1008 3234
rect 1550 3214 1554 3223
rect 1569 3214 1573 3270
rect 1850 3261 2009 3266
rect 1812 3241 1817 3247
rect 1741 3234 1744 3238
rect 2005 3235 2009 3261
rect 1550 3210 1573 3214
rect 1703 3231 1744 3234
rect 1995 3231 2009 3235
rect 1550 3208 1554 3210
rect 1688 3177 1692 3185
rect 1703 3177 1707 3231
rect 2175 3180 2179 3188
rect 2264 3180 2269 3295
rect 1629 3171 1632 3175
rect 1605 3168 1632 3171
rect 1688 3173 1707 3177
rect 2116 3174 2119 3178
rect 1688 3170 1692 3173
rect 2060 3171 2119 3174
rect 2175 3176 2269 3180
rect 2175 3173 2179 3176
rect 1416 3149 1524 3153
rect 1162 3140 1165 3144
rect 1137 3137 1165 3140
rect 483 3127 665 3132
rect 483 2785 489 3127
rect 661 3082 665 3127
rect 949 3129 1008 3133
rect 1047 3130 1050 3134
rect 949 3099 953 3129
rect 939 3095 953 3099
rect 769 3089 774 3094
rect 691 3082 694 3086
rect 661 3079 694 3082
rect 1003 3051 1008 3129
rect 1015 3127 1050 3130
rect 1015 3107 1021 3127
rect 1015 3100 1021 3102
rect 1137 3069 1145 3137
rect 1416 3102 1422 3149
rect 1520 3122 1524 3149
rect 1605 3137 1610 3168
rect 1605 3133 2008 3137
rect 1509 3118 1524 3122
rect 1554 3118 1558 3126
rect 1605 3118 1610 3133
rect 1554 3114 1610 3118
rect 1554 3111 1558 3114
rect 2004 3107 2008 3133
rect 1994 3103 2008 3107
rect 1220 3097 1422 3102
rect 2039 3102 2043 3111
rect 2060 3102 2063 3171
rect 2039 3099 2063 3102
rect 1220 3077 1225 3097
rect 2039 3096 2043 3099
rect 1003 3044 1163 3051
rect 2149 3048 2250 3051
rect 2149 3034 2156 3048
rect 561 3027 662 3030
rect 561 3009 568 3027
rect 524 3001 568 3009
rect 524 2856 532 3001
rect 545 2982 547 2987
rect 545 2946 552 2982
rect 545 2901 552 2941
rect 561 2931 568 3001
rect 658 2992 662 3027
rect 913 3029 1014 3032
rect 913 3000 920 3029
rect 873 2994 920 3000
rect 1010 2994 1014 3029
rect 1474 3029 1575 3032
rect 1474 3000 1481 3029
rect 1431 2996 1481 3000
rect 745 2947 751 2951
rect 710 2944 748 2947
rect 655 2901 660 2926
rect 710 2928 715 2944
rect 545 2895 660 2901
rect 524 2822 532 2850
rect 628 2822 633 2895
rect 873 2842 879 2994
rect 897 2984 899 2989
rect 897 2903 904 2984
rect 913 2933 920 2994
rect 1175 2978 1264 2983
rect 1096 2949 1099 2953
rect 1062 2946 1099 2949
rect 1007 2903 1012 2928
rect 1062 2930 1067 2946
rect 1431 2936 1436 2996
rect 897 2897 1012 2903
rect 974 2889 979 2897
rect 974 2876 979 2884
rect 974 2872 1021 2876
rect 1017 2842 1021 2872
rect 873 2837 887 2842
rect 894 2837 939 2842
rect 1006 2838 1021 2842
rect 1431 2843 1436 2930
rect 1458 2903 1465 2984
rect 1474 2933 1481 2996
rect 1571 2994 1575 3029
rect 2133 3003 2135 3008
rect 1657 2949 1660 2953
rect 1735 2951 1740 2956
rect 1623 2946 1660 2949
rect 1568 2903 1573 2928
rect 1623 2930 1628 2946
rect 2133 2922 2140 3003
rect 2149 2952 2156 3025
rect 2246 3013 2250 3048
rect 2332 2968 2335 2972
rect 2298 2965 2335 2968
rect 2243 2922 2248 2947
rect 2284 2948 2288 2956
rect 2298 2948 2303 2965
rect 2284 2944 2303 2948
rect 2284 2941 2288 2944
rect 2133 2916 2248 2922
rect 1458 2897 1573 2903
rect 2236 2905 2241 2916
rect 1566 2882 1571 2897
rect 1566 2843 1571 2877
rect 2236 2873 2241 2900
rect 2226 2869 2241 2873
rect 2271 2869 2275 2877
rect 2425 2869 2429 3304
rect 2271 2865 2429 2869
rect 2271 2862 2275 2865
rect 1431 2838 1500 2843
rect 1556 2839 1571 2843
rect 524 2817 585 2822
rect 619 2818 633 2822
rect 678 2785 683 2813
rect 483 2780 683 2785
<< m3contact >>
rect 1094 3741 1099 3751
rect 2451 3895 2458 3900
rect 1867 3757 1873 3763
rect 549 3485 555 3491
rect 1812 3247 1817 3253
rect 769 3094 774 3099
rect 1015 3102 1021 3107
rect 545 2941 552 2946
rect 524 2850 532 2856
rect 1431 2930 1436 2936
rect 974 2884 979 2889
rect 887 2837 894 2842
rect 2149 3025 2156 3034
rect 1740 2951 1745 2956
rect 2236 2900 2241 2905
rect 1566 2877 1571 2882
<< metal3 >>
rect 1796 3895 2451 3900
rect 1024 3741 1094 3751
rect 512 3485 549 3491
rect 1024 3490 1035 3741
rect 1796 3738 1801 3895
rect 1796 3731 1817 3738
rect 512 3345 517 3485
rect 373 3338 517 3345
rect 512 3147 517 3338
rect 769 3483 1035 3490
rect 512 3141 614 3147
rect 609 3090 614 3141
rect 769 3099 774 3483
rect 1423 3353 1521 3358
rect 1423 3244 1428 3353
rect 1517 3325 1521 3353
rect 1506 3321 1521 3325
rect 1812 3253 1817 3731
rect 1008 3240 1428 3244
rect 1442 3246 1518 3251
rect 979 3204 983 3212
rect 1008 3204 1012 3240
rect 979 3200 1012 3204
rect 979 3197 983 3200
rect 1008 3134 1012 3200
rect 1008 3130 1040 3134
rect 1442 3107 1447 3246
rect 1513 3219 1518 3246
rect 1505 3215 1518 3219
rect 1021 3102 1447 3107
rect 600 3086 614 3090
rect 1867 2956 1873 3757
rect 1745 2951 1873 2956
rect 2079 3025 2149 3034
rect 373 2941 545 2946
rect 1425 2930 1431 2936
rect 979 2884 1111 2889
rect 373 2850 524 2856
rect 887 2690 894 2837
rect 1106 2690 1111 2884
rect 1425 2811 1430 2930
rect 1571 2877 1856 2882
rect 1851 2811 1856 2877
rect 2079 2832 2092 3025
rect 2241 2900 2628 2905
rect 2622 2832 2628 2900
<< labels >>
rlabel pdcontact 1544 2850 1548 2860 1 g2n
rlabel space 2637 3824 2641 3831 1 or1s3
rlabel metal2 2544 3309 2549 3313 1 c4
rlabel pdcontact 2537 3321 2541 3331 1 c4
rlabel ndcontact 2537 3301 2541 3306 1 c4
rlabel pdcontact 2175 3188 2179 3198 1 or2c4
rlabel ndcontact 2175 3168 2179 3173 1 or2c4
rlabel polycontact 1987 3477 1991 3481 1 p2p1g0
rlabel pdcontact 2035 3362 2039 3372 1 p3p2p1p0c0
rlabel ndcontact 2035 3342 2039 3347 1 p3p2p1p0c0
rlabel polycontact 1986 3354 1990 3358 1 p2p1p0c0
rlabel pdcontact 2039 3111 2043 3121 1 p3p2g1
rlabel ndcontact 2039 3091 2043 3096 1 p3p2g1
rlabel polycontact 1990 3103 1994 3107 1 p2g1
rlabel space 2335 2965 2339 2972 1 or1p3
rlabel pdcontact 1688 3185 1692 3195 1 or2c3
rlabel ndcontact 1688 3165 1692 3170 1 or2c3
rlabel polycontact 1502 3321 1506 3325 1 p1g0
rlabel pdcontact 1550 3223 1554 3233 1 p2p1p0c0
rlabel ndcontact 1550 3203 1554 3208 1 p2p1p0c0
rlabel polycontact 1501 3215 1505 3219 1 p1p0c0
rlabel polycontact 1660 2949 1664 2953 1 or1p2
rlabel ndcontact 2271 2857 2275 2862 1 g3
rlabel pdcontact 2271 2877 2275 2887 1 g3
rlabel polycontact 1552 2839 1556 2843 1 b2
rlabel metal1 2697 3829 2708 3833 1 s3
rlabel ndcontact 2693 3821 2697 3826 1 s3
rlabel pdcontact 2693 3841 2697 3851 1 s3
rlabel pdiffusion 2634 3838 2640 3858 1 orpms3
rlabel polycontact 2677 3829 2681 3833 1 s3n
rlabel ndcontact 2634 3813 2640 3818 1 s3n
rlabel pdcontact 2644 3838 2648 3858 1 s3n
rlabel pdcontact 2586 3815 2590 3825 1 or1s3
rlabel ndcontact 2586 3795 2590 3800 1 or1s3
rlabel polycontact 2627 3827 2631 3831 1 or2s3
rlabel ndcontact 2584 3861 2588 3866 1 or2s3
rlabel pdcontact 2584 3881 2588 3891 1 or2s3
rlabel ndiffusion 2526 3855 2532 3865 1 and1nms3
rlabel ndiffusion 2528 3789 2534 3799 1 and2nms3
rlabel polycontact 2570 3803 2574 3807 1 and2ns3
rlabel ndcontact 2538 3789 2542 3799 1 and2ns3
rlabel pdcontact 2529 3818 2533 3828 1 and2ns3
rlabel polycontact 2568 3869 2572 3873 1 and1ns3
rlabel ndcontact 2536 3855 2540 3865 1 and1ns3
rlabel pdcontact 2527 3884 2531 3894 1 and1ns3
rlabel polycontact 2519 3873 2523 3877 1 p3not
rlabel pdcontact 2490 3874 2494 3884 1 p3not
rlabel ndcontact 2490 3854 2494 3859 1 p3not
rlabel polycontact 2521 3807 2525 3811 1 c3not
rlabel pdcontact 2490 3818 2494 3828 1 c3not
rlabel ndcontact 2490 3798 2494 3803 1 c3not
rlabel polycontact 2535 3873 2539 3877 1 c3
rlabel polycontact 2474 3806 2478 3810 1 c3
rlabel polycontact 2537 3807 2541 3811 1 p3
rlabel polycontact 2474 3862 2478 3866 1 p3
rlabel metal1 2075 3811 2086 3815 1 s2
rlabel pdcontact 2071 3823 2075 3833 1 s2
rlabel ndcontact 2071 3803 2075 3808 1 s2
rlabel polycontact 2055 3811 2059 3815 1 s2n
rlabel ndcontact 2012 3795 2018 3800 1 s2n
rlabel pdcontact 2022 3820 2026 3840 1 s2n
rlabel pdiffusion 2012 3820 2018 3840 1 orpms2
rlabel polycontact 2015 3809 2019 3813 1 or1s2
rlabel pdcontact 1964 3797 1968 3807 1 or1s2
rlabel ndcontact 1964 3777 1968 3782 1 or1s2
rlabel polycontact 2005 3809 2009 3813 1 or2s2
rlabel ndcontact 1962 3843 1966 3848 1 or2s2
rlabel pdcontact 1962 3863 1966 3873 1 or2s2
rlabel polycontact 1948 3785 1952 3789 1 and2ns2
rlabel ndiffusion 1906 3771 1912 3781 1 and2nms2
rlabel ndcontact 1916 3771 1920 3781 1 and2ns2
rlabel pdcontact 1907 3800 1911 3810 1 and2ns2
rlabel polycontact 1946 3851 1950 3855 1 and1ns2
rlabel ndcontact 1914 3837 1918 3847 1 and1ns2
rlabel ndiffusion 1904 3837 1910 3847 1 and1nms2
rlabel pdcontact 1905 3866 1909 3876 1 and1ns2
rlabel polycontact 1897 3855 1901 3859 1 p2not
rlabel pdcontact 1868 3856 1872 3866 1 p2not
rlabel ndcontact 1868 3836 1872 3841 1 p2not
rlabel polycontact 1913 3855 1917 3859 1 c2
rlabel polycontact 1852 3844 1856 3848 1 p2
rlabel polycontact 1915 3789 1919 3793 1 p2
rlabel polycontact 1899 3789 1903 3793 1 c2not
rlabel pdcontact 1868 3800 1872 3810 1 c2not
rlabel ndcontact 1868 3780 1872 3785 1 c2not
rlabel polycontact 1852 3788 1856 3792 1 c2
rlabel pdcontact 2022 3239 2026 3249 1 vdd
rlabel polycontact 1668 3275 1672 3279 1 orc3n
rlabel metal1 1642 3267 1652 3271 1 orc3n
rlabel ndcontact 1625 3259 1631 3264 1 orc3n
rlabel pdcontact 1635 3284 1639 3304 1 orc3n
rlabel pdcontact 1639 3182 1643 3202 1 or2c3n
rlabel ndcontact 1629 3157 1635 3162 1 or2c3n
rlabel metal1 1643 3165 1652 3169 1 or2c3n
rlabel polycontact 1672 3173 1676 3177 1 or2c3n
rlabel metal2 1694 3173 1703 3177 1 or2c3
rlabel polycontact 1744 3234 1748 3238 1 or2c3
rlabel polycontact 1734 3234 1738 3238 1 orc3
rlabel metal1 1691 3275 1701 3279 1 orc3
rlabel ndcontact 1684 3267 1688 3272 1 orc3
rlabel pdcontact 1684 3287 1688 3297 1 orc3
rlabel ndcontact 2519 3301 2523 3306 1 gnd
rlabel ndcontact 2488 3293 2492 3298 1 gnd
rlabel ndcontact 2470 3293 2474 3298 1 gnd
rlabel pdcontact 2519 3321 2523 3331 1 vdd
rlabel pdcontact 2470 3318 2474 3338 1 vdd
rlabel polycontact 2521 3309 2525 3313 1 coutn
rlabel metal1 2493 3301 2498 3305 1 coutn
rlabel ndcontact 2478 3293 2484 3298 1 coutn
rlabel pdcontact 2488 3318 2492 3338 1 coutn
rlabel pdiffusion 2478 3318 2484 3338 1 or0pmc4
rlabel polycontact 2471 3307 2475 3311 1 or1c4
rlabel metal1 2362 3300 2370 3304 1 or1c4
rlabel ndcontact 2352 3292 2356 3297 1 or1c4
rlabel pdcontact 2352 3312 2356 3322 1 or1c4
rlabel polycontact 2336 3300 2340 3304 1 or1c4n
rlabel metal1 2314 3292 2318 3296 1 or1c4n
rlabel ndcontact 2293 3284 2299 3289 1 or1c4n
rlabel pdcontact 2303 3309 2307 3329 1 or1c4n
rlabel ndcontact 2334 3292 2338 3297 1 gnd
rlabel ndcontact 2303 3284 2307 3289 1 gnd
rlabel ndcontact 2285 3284 2289 3289 1 gnd
rlabel pdcontact 2334 3312 2338 3322 1 vdd
rlabel pdcontact 2285 3309 2289 3329 1 vdd
rlabel pdiffusion 2293 3309 2299 3329 1 or1pmc4
rlabel polycontact 2296 3298 2300 3302 1 or2c4
rlabel metal2 2199 3176 2207 3180 1 or2c4
rlabel polycontact 2159 3176 2163 3180 1 or2c4n
rlabel metal1 2133 3168 2139 3172 1 or2c4n
rlabel ndcontact 2116 3160 2122 3165 1 or2c4n
rlabel pdcontact 2126 3185 2130 3205 1 or2c4n
rlabel pdiffusion 2116 3185 2122 3205 1 or2pmc4
rlabel ndcontact 2157 3168 2161 3173 1 gnd
rlabel ndcontact 2126 3160 2130 3165 1 gnd
rlabel ndcontact 2108 3160 2112 3165 1 gnd
rlabel pdcontact 2157 3188 2161 3198 1 vdd
rlabel pdcontact 2108 3185 2112 3205 1 vdd
rlabel polycontact 2286 3298 2290 3302 1 or3c4
rlabel metal1 2185 3420 2190 3424 1 or3c4
rlabel ndcontact 2176 3412 2180 3417 1 or3c4
rlabel pdcontact 2176 3432 2180 3442 1 or3c4
rlabel polycontact 2160 3420 2164 3424 1 or3nc4
rlabel metal1 2140 3412 2144 3420 1 or3nc4
rlabel ndcontact 2117 3404 2123 3409 1 or3nc4
rlabel pdcontact 2127 3429 2131 3449 1 or3nc4
rlabel pdiffusion 2117 3429 2123 3449 1 or3pmc4
rlabel ndcontact 2158 3412 2162 3417 1 gnd
rlabel ndcontact 2127 3404 2131 3409 1 gnd
rlabel ndcontact 2109 3404 2113 3409 1 gnd
rlabel pdcontact 2158 3432 2162 3442 1 vdd
rlabel pdcontact 2109 3429 2113 3449 1 vdd
rlabel polycontact 2110 3418 2114 3422 1 p3p2p1g0
rlabel ndcontact 2022 3219 2026 3224 1 gnd
rlabel pdcontact 2021 3111 2025 3121 1 vdd
rlabel ndcontact 2021 3091 2025 3096 1 gnd
rlabel ndcontact 1973 3085 1977 3095 1 gnd
rlabel pdcontact 1991 3114 1995 3124 1 vdd
rlabel pdcontact 1973 3114 1977 3124 1 vdd
rlabel polycontact 1971 3476 1975 3481 1 p3
rlabel metal1 2049 3473 2059 3477 1 p3p2p1g0
rlabel pdcontact 2036 3485 2040 3495 1 p3p2p1g0
rlabel ndcontact 2036 3465 2040 3470 1 p3p2p1g0
rlabel ndcontact 2018 3465 2022 3470 1 gnd
rlabel ndiffusion 1978 3459 1984 3469 1 and4nmc4
rlabel polycontact 2020 3473 2024 3477 1 p3p2p1g0n
rlabel metal1 1994 3469 2004 3473 1 p3p2p1g0n
rlabel ndcontact 1988 3459 1992 3469 1 p3p2p1g0n
rlabel pdcontact 1979 3488 1983 3498 1 p3p2p1g0n
rlabel pdcontact 2018 3485 2022 3495 1 vdd
rlabel pdcontact 1988 3488 1992 3498 1 vdd
rlabel pdcontact 1970 3488 1974 3498 1 vdd
rlabel ndcontact 1970 3459 1974 3469 1 gnd
rlabel ndcontact 1969 3336 1973 3346 1 gnd
rlabel ndcontact 2017 3342 2021 3347 1 gnd
rlabel polycontact 2120 3418 2124 3422 1 p3p2p1p0c0
rlabel metal2 2045 3350 2056 3353 1 p3p2p1p0c0
rlabel polycontact 2019 3350 2023 3354 1 p3p2p1p0c0n
rlabel ndiffusion 1977 3336 1983 3346 1 and3nmc4
rlabel ndcontact 1987 3336 1991 3346 1 p3p2p1p0c0n
rlabel pdcontact 1978 3365 1982 3375 1 p3p2p1p0c0n
rlabel pdcontact 1987 3365 1991 3375 1 vdd
rlabel pdcontact 1969 3365 1973 3375 1 vdd
rlabel pdcontact 2017 3362 2021 3372 1 vdd
rlabel polycontact 2109 3174 2113 3178 1 p3g2
rlabel metal1 2053 3227 2060 3231 1 p3g2
rlabel ndcontact 2040 3219 2044 3224 1 p3g2
rlabel pdcontact 2040 3239 2044 3249 1 p3g2
rlabel polycontact 2024 3227 2028 3231 1 p3g2n
rlabel metal1 2000 3223 2008 3227 1 p3g2n
rlabel ndcontact 1992 3213 1996 3223 1 p3g2n
rlabel pdcontact 1983 3242 1987 3252 1 p3g2n
rlabel pdcontact 1992 3242 1996 3252 1 vdd
rlabel pdcontact 1974 3242 1978 3252 1 vdd
rlabel ndcontact 1974 3213 1978 3223 1 gnd
rlabel ndiffusion 1982 3213 1988 3223 1 and2nmc4
rlabel ndiffusion 1981 3085 1987 3095 1 and1nmc4
rlabel metal2 2051 3099 2060 3102 1 p2p3g1
rlabel polycontact 2023 3099 2027 3103 1 p2p3g1n
rlabel ndcontact 1991 3085 1995 3095 1 p2p3g1n
rlabel pdcontact 1982 3114 1986 3124 1 p2p3g1n
rlabel polycontact 2481 3307 2485 3311 1 g3
rlabel polycontact 1970 3354 1974 3358 1 p3
rlabel polycontact 1975 3231 1979 3235 1 p3
rlabel polycontact 1974 3103 1978 3107 1 p3
rlabel metal1 1807 3236 1812 3240 1 c3
rlabel ndcontact 1800 3228 1804 3233 1 c3
rlabel pdcontact 1800 3248 1804 3258 1 c3
rlabel polycontact 1784 3236 1788 3240 1 c3n
rlabel metal1 1764 3228 1768 3240 1 c3n
rlabel ndcontact 1741 3220 1747 3225 1 c3n
rlabel pdcontact 1751 3245 1755 3265 1 c3n
rlabel pdiffusion 1741 3245 1747 3265 1 or1pmc3
rlabel pdiffusion 1629 3182 1635 3202 1 or2pmc3
rlabel polycontact 1632 3171 1636 3175 1 p2g1
rlabel polycontact 1622 3171 1626 3175 1 g2
rlabel pdiffusion 1625 3284 1631 3304 1 or3pmc3
rlabel polycontact 1618 3273 1622 3277 1 p2p1g0
rlabel polycontact 1628 3273 1632 3277 1 p2p1p0c0
rlabel ndiffusion 1493 3303 1499 3313 1 and3nmc3
rlabel metal1 1555 3317 1567 3321 1 p2p1g0
rlabel ndcontact 1551 3309 1555 3314 1 p2p1g0
rlabel pdcontact 1551 3329 1555 3339 1 p2p1g0
rlabel polycontact 1535 3317 1539 3321 1 p2p1g0n
rlabel ndcontact 1503 3303 1507 3313 1 p2p1g0n
rlabel pdcontact 1494 3332 1498 3342 1 p2p1g0n
rlabel metal2 1558 3114 1569 3118 1 p2g1
rlabel polycontact 1538 3114 1542 3118 1 p2g1n
rlabel metal1 1514 3110 1522 3114 1 p2g1n
rlabel ndcontact 1506 3100 1510 3110 1 p2g1n
rlabel pdcontact 1497 3129 1501 3139 1 p2g1n
rlabel ndiffusion 1496 3100 1502 3110 1 and1nmc3
rlabel ndiffusion 1492 3197 1498 3207 1 and2nmc3
rlabel metal2 1556 3210 1566 3214 1 p2p1p0c0
rlabel polycontact 1534 3211 1538 3215 1 p2p1p0c0n
rlabel ndcontact 1502 3197 1506 3207 1 p2p1p0c0n
rlabel pdcontact 1493 3226 1497 3236 1 p2p1p0c0n
rlabel polycontact 1486 3321 1490 3325 1 p2
rlabel polycontact 1485 3215 1489 3219 1 p2
rlabel polycontact 1489 3118 1493 3122 1 p2
rlabel metal2 2278 2865 2295 2869 1 g3
rlabel ndiffusion 2213 2851 2219 2861 1 and1nmg3
rlabel polycontact 2255 2865 2259 2869 1 g3n
rlabel ndcontact 2223 2851 2227 2861 1 g3n
rlabel pdcontact 2214 2880 2218 2890 1 g3n
rlabel polycontact 2206 2869 2210 2873 1 a3
rlabel metal1 1608 2835 1623 2839 1 g2
rlabel pdcontact 1601 2847 1605 2857 1 g2
rlabel ndcontact 1601 2827 1605 2832 1 g2
rlabel ndiffusion 1543 2821 1549 2831 1 and1nmg2
rlabel polycontact 1585 2835 1589 2839 1 g2n
rlabel ndcontact 1553 2821 1557 2831 1 g2n
rlabel polycontact 1536 2838 1540 2843 1 a2
rlabel ndcontact 1583 2827 1587 2832 1 gnd
rlabel ndcontact 1535 2821 1539 2831 1 gnd
rlabel ndcontact 2205 2851 2209 2861 1 gnd
rlabel ndcontact 2253 2857 2257 2862 1 gnd
rlabel metal1 2247 2848 2281 2851 1 gnd
rlabel metal1 2199 2844 2233 2847 1 gnd
rlabel metal1 1577 2818 1611 2821 1 gnd
rlabel metal1 1529 2814 1563 2817 1 gnd
rlabel metal1 1577 2863 1611 2867 1 vdd
rlabel metal1 1529 2865 1563 2869 1 vdd
rlabel metal1 2199 2895 2233 2899 1 vdd
rlabel metal1 2247 2893 2281 2897 1 vdd
rlabel pdcontact 2253 2877 2257 2887 1 vdd
rlabel pdcontact 2223 2880 2227 2890 1 vdd
rlabel pdcontact 2205 2880 2209 2890 1 vdd
rlabel pdcontact 1583 2847 1587 2857 1 vdd
rlabel pdcontact 1553 2850 1557 2860 1 vdd
rlabel pdcontact 1535 2850 1539 2860 1 vdd
rlabel pdcontact 1533 3329 1537 3339 1 vdd
rlabel pdcontact 1503 3332 1507 3342 1 vdd
rlabel pdcontact 1485 3332 1489 3342 1 vdd
rlabel pdcontact 1502 3226 1506 3236 1 vdd
rlabel pdcontact 1484 3226 1488 3236 1 vdd
rlabel pdcontact 1506 3129 1510 3139 1 vdd
rlabel pdcontact 1488 3129 1492 3139 1 vdd
rlabel pdcontact 1536 3126 1540 3136 1 vdd
rlabel pdcontact 1532 3223 1536 3233 1 vdd
rlabel pdcontact 1670 3185 1674 3195 1 vdd
rlabel pdcontact 1666 3287 1670 3297 1 vdd
rlabel pdcontact 1617 3284 1621 3304 1 vdd
rlabel pdcontact 1621 3182 1625 3202 1 vdd
rlabel pdcontact 1733 3245 1737 3265 1 vdd
rlabel pdcontact 1782 3248 1786 3258 1 vdd
rlabel ndcontact 1782 3228 1786 3233 1 gnd
rlabel ndcontact 1751 3220 1755 3225 1 gnd
rlabel ndcontact 1733 3220 1737 3225 1 gnd
rlabel ndcontact 1670 3165 1674 3170 1 gnd
rlabel ndcontact 1666 3267 1670 3272 1 gnd
rlabel ndcontact 1635 3259 1639 3264 1 gnd
rlabel ndcontact 1617 3259 1621 3264 1 gnd
rlabel ndcontact 1639 3157 1643 3162 1 gnd
rlabel ndcontact 1621 3157 1625 3162 1 gnd
rlabel ndcontact 1536 3106 1540 3111 1 gnd
rlabel ndcontact 1532 3203 1536 3208 1 gnd
rlabel ndcontact 1533 3309 1537 3314 1 gnd
rlabel ndcontact 1485 3303 1489 3313 1 gnd
rlabel ndcontact 1484 3197 1488 3207 1 gnd
rlabel ndcontact 1488 3100 1492 3110 1 gnd
rlabel metal1 1530 3097 1564 3100 1 gnd
rlabel metal1 1482 3093 1516 3096 1 gnd
rlabel metal1 1527 3300 1561 3303 1 gnd
rlabel metal1 1479 3296 1513 3299 1 gnd
rlabel metal1 1478 3190 1512 3193 1 gnd
rlabel metal1 1526 3194 1560 3197 1 gnd
rlabel metal1 1664 3156 1698 3159 1 gnd
rlabel metal1 1615 3148 1649 3151 1 gnd
rlabel metal1 1660 3258 1694 3261 1 gnd
rlabel metal1 1611 3250 1645 3253 1 gnd
rlabel metal1 1727 3211 1761 3214 1 gnd
rlabel metal1 1776 3219 1810 3222 1 gnd
rlabel metal1 2015 3082 2049 3085 1 gnd
rlabel metal1 1967 3078 2001 3081 1 gnd
rlabel metal1 2016 3210 2050 3213 1 gnd
rlabel metal1 1968 3206 2002 3209 1 gnd
rlabel metal1 2011 3333 2045 3336 1 gnd
rlabel metal1 1963 3329 1997 3332 1 gnd
rlabel metal1 2012 3456 2046 3459 1 gnd
rlabel metal1 1964 3452 1998 3455 1 gnd
rlabel metal1 2152 3403 2186 3406 1 gnd
rlabel metal1 2103 3395 2137 3398 1 gnd
rlabel metal1 2151 3159 2185 3162 1 gnd
rlabel metal1 2102 3151 2136 3154 1 gnd
rlabel metal1 2279 3275 2313 3278 1 gnd
rlabel metal1 2328 3283 2362 3286 1 gnd
rlabel metal1 2464 3284 2498 3287 1 gnd
rlabel metal1 2513 3292 2547 3295 1 gnd
rlabel metal1 2513 3337 2547 3341 1 vdd
rlabel metal1 2464 3346 2498 3350 1 vdd
rlabel metal1 2328 3328 2362 3332 1 vdd
rlabel metal1 2279 3337 2313 3341 1 vdd
rlabel metal1 2152 3448 2186 3452 1 vdd
rlabel metal1 2103 3457 2137 3461 1 vdd
rlabel metal1 2012 3501 2046 3505 1 vdd
rlabel metal1 1964 3503 1998 3507 1 vdd
rlabel metal1 2011 3378 2045 3382 1 vdd
rlabel metal1 1963 3380 1997 3384 1 vdd
rlabel metal1 2151 3204 2185 3208 1 vdd
rlabel metal1 2102 3213 2136 3217 1 vdd
rlabel metal1 2015 3127 2049 3131 1 vdd
rlabel metal1 1967 3129 2001 3133 1 vdd
rlabel metal1 2016 3255 2050 3259 1 vdd
rlabel metal1 1968 3257 2002 3261 1 vdd
rlabel metal1 1776 3264 1810 3268 1 vdd
rlabel metal1 1727 3273 1761 3277 1 vdd
rlabel metal1 1664 3201 1698 3205 1 vdd
rlabel metal1 1615 3210 1649 3214 1 vdd
rlabel metal1 1660 3303 1694 3307 1 vdd
rlabel metal1 1611 3312 1645 3316 1 vdd
rlabel metal1 1530 3142 1564 3146 1 vdd
rlabel metal1 1482 3144 1516 3148 1 vdd
rlabel metal1 1526 3239 1560 3243 1 vdd
rlabel metal1 1478 3241 1512 3245 1 vdd
rlabel metal1 1527 3345 1561 3349 1 vdd
rlabel metal1 1479 3347 1513 3351 1 vdd
rlabel metal1 2395 2970 2406 2974 1 p3
rlabel pdcontact 2391 2982 2395 2992 1 p3
rlabel ndcontact 2391 2962 2395 2967 1 p3
rlabel polycontact 2375 2970 2379 2974 1 outnp3
rlabel pdcontact 2342 2979 2346 2999 1 outnp3
rlabel ndcontact 2332 2954 2338 2959 1 outnp3
rlabel pdiffusion 2332 2979 2338 2999 1 orpmp3
rlabel ndcontact 2284 2936 2288 2941 1 or1p3
rlabel pdcontact 2284 2956 2288 2966 1 or1p3
rlabel ndcontact 2282 3002 2286 3007 1 or2p3
rlabel pdcontact 2282 3022 2286 3032 1 or2p3
rlabel polycontact 2235 2948 2239 2952 1 b3
rlabel ndiffusion 2226 2930 2232 2940 1 and2nmp3
rlabel polycontact 2268 2944 2272 2948 1 and2np3
rlabel ndcontact 2236 2930 2240 2940 1 and2np3
rlabel pdcontact 2227 2959 2231 2969 1 and2np3
rlabel ndiffusion 2224 2996 2230 3006 1 and1nmp3
rlabel polycontact 2233 3014 2237 3018 1 a3
rlabel polycontact 2266 3010 2270 3014 1 and1np3
rlabel ndcontact 2234 2996 2238 3006 1 and1np3
rlabel pdcontact 2225 3025 2229 3035 1 and1np3
rlabel polycontact 2219 2948 2223 2952 1 a3not
rlabel pdcontact 2188 2959 2192 2969 1 a3not
rlabel ndcontact 2188 2939 2192 2944 1 a3not
rlabel polycontact 2172 2947 2176 2951 1 a3
rlabel polycontact 2217 3014 2221 3018 1 b3not
rlabel pdcontact 2188 3015 2192 3025 1 b3not
rlabel ndcontact 2188 2995 2192 3000 1 b3not
rlabel polycontact 2172 3003 2176 3007 1 b3
rlabel metal1 1720 2951 1730 2955 1 p2
rlabel pdcontact 1716 2963 1720 2973 1 p2
rlabel ndcontact 1716 2943 1720 2948 1 p2
rlabel polycontact 1700 2951 1704 2955 1 outnp2
rlabel pdcontact 1667 2960 1671 2980 1 outnp2
rlabel ndcontact 1657 2935 1663 2940 1 outnp2
rlabel pdiffusion 1657 2960 1663 2980 1 orpmp2
rlabel ndcontact 1609 2917 1613 2922 1 or1p2
rlabel pdcontact 1609 2937 1613 2947 1 or1p2
rlabel polycontact 1650 2949 1654 2953 1 or2p2
rlabel ndcontact 1607 2983 1611 2988 1 or2p2
rlabel pdcontact 1607 3003 1611 3013 1 or2p2
rlabel ndiffusion 1549 2977 1555 2987 1 and1nmp2
rlabel polycontact 1558 2995 1562 2999 1 a2
rlabel polycontact 1591 2991 1595 2995 1 and1np2
rlabel ndcontact 1559 2977 1563 2987 1 and1np2
rlabel pdcontact 1550 3006 1554 3016 1 and1np2
rlabel polycontact 1542 2995 1546 2999 1 b2not
rlabel pdcontact 1513 2996 1517 3006 1 b2not
rlabel ndcontact 1513 2976 1517 2981 1 b2not
rlabel polycontact 1497 2984 1501 2989 1 b2
rlabel ndiffusion 1551 2911 1557 2921 1 and2nmp2
rlabel polycontact 1593 2925 1597 2929 1 and2np2
rlabel ndcontact 1561 2911 1565 2921 1 and2np2
rlabel polycontact 1560 2929 1564 2933 1 b2
rlabel pdcontact 1552 2940 1556 2950 1 and2np2
rlabel polycontact 1544 2929 1548 2933 1 a2not
rlabel pdcontact 1513 2940 1517 2950 1 a2not
rlabel ndcontact 1513 2920 1517 2925 1 a2not
rlabel polycontact 1497 2928 1501 2932 1 a2
rlabel ndcontact 2566 3861 2570 3866 1 gnd
rlabel metal1 2560 3852 2594 3855 1 gnd
rlabel metal1 2514 3782 2545 3785 1 gnd
rlabel ndcontact 2518 3855 2522 3865 1 gnd
rlabel ndcontact 2472 3854 2476 3859 1 gnd
rlabel metal1 2512 3848 2546 3851 1 gnd
rlabel metal1 2466 3845 2500 3848 1 gnd
rlabel metal1 2466 3789 2500 3792 1 gnd
rlabel ndcontact 2472 3798 2476 3803 1 gnd
rlabel ndcontact 2568 3795 2572 3800 1 gnd
rlabel ndcontact 2520 3789 2524 3799 1 gnd
rlabel metal1 2562 3786 2596 3789 1 gnd
rlabel metal1 2669 3812 2703 3815 1 gnd
rlabel ndcontact 2675 3821 2679 3826 1 gnd
rlabel ndcontact 2644 3813 2648 3818 1 gnd
rlabel ndcontact 2626 3813 2630 3818 1 gnd
rlabel metal1 2620 3804 2654 3807 1 gnd
rlabel pdcontact 2675 3841 2679 3851 1 vdd
rlabel metal1 2669 3857 2703 3861 1 vdd
rlabel pdcontact 2626 3838 2630 3858 1 vdd
rlabel metal1 2620 3866 2654 3870 1 vdd
rlabel pdcontact 2568 3815 2572 3825 1 vdd
rlabel metal1 2562 3831 2596 3835 1 vdd
rlabel pdcontact 2538 3818 2542 3828 1 vdd
rlabel pdcontact 2520 3818 2524 3828 1 vdd
rlabel metal1 2514 3833 2548 3837 1 vdd
rlabel pdcontact 2472 3818 2476 3828 1 vdd
rlabel metal1 2466 3834 2500 3838 1 vdd
rlabel pdcontact 2566 3881 2570 3891 1 vdd
rlabel metal1 2560 3897 2594 3901 5 vdd
rlabel pdcontact 2536 3884 2540 3894 1 vdd
rlabel pdcontact 2518 3884 2522 3894 1 vdd
rlabel metal1 2512 3899 2546 3903 5 vdd
rlabel pdcontact 2472 3874 2476 3884 1 vdd
rlabel metal1 2466 3890 2500 3894 1 vdd
rlabel ndcontact 1944 3843 1948 3848 1 gnd
rlabel metal1 1938 3834 1972 3837 1 gnd
rlabel metal1 1892 3764 1923 3767 1 gnd
rlabel ndcontact 1896 3837 1900 3847 1 gnd
rlabel ndcontact 1850 3836 1854 3841 1 gnd
rlabel metal1 1890 3830 1924 3833 1 gnd
rlabel metal1 1844 3827 1878 3830 1 gnd
rlabel metal1 1844 3771 1878 3774 1 gnd
rlabel ndcontact 1850 3780 1854 3785 1 gnd
rlabel ndcontact 1946 3777 1950 3782 1 gnd
rlabel ndcontact 1898 3771 1902 3781 1 gnd
rlabel metal1 1940 3768 1974 3771 1 gnd
rlabel metal1 2047 3794 2081 3797 1 gnd
rlabel ndcontact 2053 3803 2057 3808 1 gnd
rlabel ndcontact 2022 3795 2026 3800 1 gnd
rlabel ndcontact 2004 3795 2008 3800 1 gnd
rlabel metal1 1998 3786 2032 3789 1 gnd
rlabel pdcontact 2053 3823 2057 3833 1 vdd
rlabel metal1 2047 3839 2081 3843 1 vdd
rlabel pdcontact 2004 3820 2008 3840 1 vdd
rlabel metal1 1998 3848 2032 3852 1 vdd
rlabel pdcontact 1946 3797 1950 3807 1 vdd
rlabel metal1 1940 3813 1974 3817 1 vdd
rlabel pdcontact 1916 3800 1920 3810 1 vdd
rlabel pdcontact 1898 3800 1902 3810 1 vdd
rlabel metal1 1892 3815 1926 3819 1 vdd
rlabel pdcontact 1850 3800 1854 3810 1 vdd
rlabel metal1 1844 3816 1878 3820 1 vdd
rlabel pdcontact 1944 3863 1948 3873 1 vdd
rlabel metal1 1938 3879 1972 3883 5 vdd
rlabel pdcontact 1914 3866 1918 3876 1 vdd
rlabel pdcontact 1896 3866 1900 3876 1 vdd
rlabel metal1 1890 3881 1924 3885 5 vdd
rlabel pdcontact 1850 3856 1854 3866 1 vdd
rlabel metal1 1844 3872 1878 3876 1 vdd
rlabel ndcontact 2264 3002 2268 3007 1 gnd
rlabel metal1 2258 2993 2292 2996 1 gnd
rlabel metal1 2212 2923 2243 2926 1 gnd
rlabel ndcontact 2216 2996 2220 3006 1 gnd
rlabel ndcontact 2170 2995 2174 3000 1 gnd
rlabel metal1 2210 2989 2244 2992 1 gnd
rlabel metal1 2164 2986 2198 2989 1 gnd
rlabel metal1 2164 2930 2198 2933 1 gnd
rlabel ndcontact 2170 2939 2174 2944 1 gnd
rlabel ndcontact 2266 2936 2270 2941 1 gnd
rlabel ndcontact 2218 2930 2222 2940 1 gnd
rlabel metal1 2260 2927 2294 2930 1 gnd
rlabel metal1 2367 2953 2401 2956 1 gnd
rlabel ndcontact 2373 2962 2377 2967 1 gnd
rlabel ndcontact 2342 2954 2346 2959 1 gnd
rlabel ndcontact 2324 2954 2328 2959 1 gnd
rlabel metal1 2318 2945 2352 2948 1 gnd
rlabel pdcontact 2373 2982 2377 2992 1 vdd
rlabel metal1 2367 2998 2401 3002 1 vdd
rlabel pdcontact 2324 2979 2328 2999 1 vdd
rlabel metal1 2318 3007 2352 3011 1 vdd
rlabel pdcontact 2266 2956 2270 2966 1 vdd
rlabel metal1 2260 2972 2294 2976 1 vdd
rlabel pdcontact 2236 2959 2240 2969 1 vdd
rlabel pdcontact 2218 2959 2222 2969 1 vdd
rlabel metal1 2212 2974 2246 2978 1 vdd
rlabel pdcontact 2170 2959 2174 2969 1 vdd
rlabel metal1 2164 2975 2198 2979 1 vdd
rlabel pdcontact 2264 3022 2268 3032 1 vdd
rlabel metal1 2258 3038 2292 3042 5 vdd
rlabel pdcontact 2234 3025 2238 3035 1 vdd
rlabel pdcontact 2216 3025 2220 3035 1 vdd
rlabel metal1 2210 3040 2244 3044 5 vdd
rlabel pdcontact 2170 3015 2174 3025 1 vdd
rlabel metal1 2164 3031 2198 3035 1 vdd
rlabel ndcontact 1589 2983 1593 2988 1 gnd
rlabel metal1 1583 2974 1617 2977 1 gnd
rlabel metal1 1537 2904 1568 2907 1 gnd
rlabel ndcontact 1541 2977 1545 2987 1 gnd
rlabel ndcontact 1495 2976 1499 2981 1 gnd
rlabel metal1 1535 2970 1569 2973 1 gnd
rlabel metal1 1489 2967 1523 2970 1 gnd
rlabel metal1 1489 2911 1523 2914 1 gnd
rlabel ndcontact 1495 2920 1499 2925 1 gnd
rlabel ndcontact 1591 2917 1595 2922 1 gnd
rlabel ndcontact 1543 2911 1547 2921 1 gnd
rlabel metal1 1585 2908 1619 2911 1 gnd
rlabel metal1 1692 2934 1726 2937 1 gnd
rlabel ndcontact 1698 2943 1702 2948 1 gnd
rlabel ndcontact 1667 2935 1671 2940 1 gnd
rlabel ndcontact 1649 2935 1653 2940 1 gnd
rlabel metal1 1643 2926 1677 2929 1 gnd
rlabel pdcontact 1698 2963 1702 2973 1 vdd
rlabel metal1 1692 2979 1726 2983 1 vdd
rlabel pdcontact 1649 2960 1653 2980 1 vdd
rlabel metal1 1643 2988 1677 2992 1 vdd
rlabel pdcontact 1591 2937 1595 2947 1 vdd
rlabel metal1 1585 2953 1619 2957 1 vdd
rlabel pdcontact 1561 2940 1565 2950 1 vdd
rlabel pdcontact 1543 2940 1547 2950 1 vdd
rlabel metal1 1537 2955 1571 2959 1 vdd
rlabel pdcontact 1495 2940 1499 2950 1 vdd
rlabel metal1 1489 2956 1523 2960 1 vdd
rlabel pdcontact 1589 3003 1593 3013 1 vdd
rlabel metal1 1583 3019 1617 3023 5 vdd
rlabel pdcontact 1559 3006 1563 3016 1 vdd
rlabel pdcontact 1541 3006 1545 3016 1 vdd
rlabel metal1 1535 3021 1569 3025 5 vdd
rlabel pdcontact 1495 2996 1499 3006 1 vdd
rlabel metal1 1489 3012 1523 3016 1 vdd
rlabel polycontact 1040 3130 1044 3134 1 p1g0
rlabel polycontact 615 2818 619 2822 1 b0
rlabel polycontact 1192 3829 1196 3833 1 p1
rlabel polycontact 586 3572 590 3576 1 c0
rlabel polycontact 649 3517 653 3521 1 c0
rlabel polycontact 963 3200 967 3204 1 p1g0n
rlabel pdcontact 979 3212 983 3222 1 p1g0
rlabel ndcontact 979 3192 983 3197 1 p1g0
rlabel polycontact 935 3095 939 3099 1 p1
rlabel polycontact 930 3204 934 3208 1 p1
rlabel metal1 1354 3785 1365 3789 1 s1
rlabel ndcontact 1350 3777 1354 3782 1 s1
rlabel pdcontact 1350 3797 1354 3807 1 s1
rlabel polycontact 1334 3785 1338 3789 1 s1n
rlabel ndcontact 1291 3769 1297 3774 1 s1n
rlabel pdcontact 1301 3794 1305 3814 1 s1n
rlabel pdiffusion 1291 3794 1297 3814 1 orpms1
rlabel pdcontact 1241 3837 1245 3847 1 or2s1
rlabel ndcontact 1241 3817 1245 3822 1 or2s1
rlabel polycontact 1294 3783 1298 3787 1 or1s1
rlabel polycontact 1284 3783 1288 3787 1 or2s1
rlabel ndcontact 1243 3751 1247 3756 1 or1s1
rlabel pdcontact 1243 3771 1247 3781 1 or1s1
rlabel ndiffusion 1185 3745 1191 3755 1 and2nms1
rlabel ndiffusion 1183 3811 1189 3821 1 and1nms1
rlabel polycontact 1225 3825 1229 3829 1 and1ns1
rlabel polycontact 1227 3759 1231 3763 1 and2ns1
rlabel ndcontact 1195 3745 1199 3755 1 and2ns1
rlabel ndcontact 1193 3811 1197 3821 1 and1ns1
rlabel pdcontact 1184 3840 1188 3850 1 and1ns1
rlabel pdcontact 1186 3774 1190 3784 1 and2ns1
rlabel polycontact 1194 3763 1198 3767 1 c1
rlabel polycontact 1178 3763 1182 3767 1 p1not
rlabel pdcontact 1147 3774 1151 3784 1 p1not
rlabel ndcontact 1147 3754 1151 3759 1 p1not
rlabel polycontact 1176 3829 1180 3833 1 c1not
rlabel pdcontact 1147 3830 1151 3840 1 c1not
rlabel ndcontact 1147 3810 1151 3815 1 c1not
rlabel polycontact 1131 3818 1135 3822 1 c1
rlabel polycontact 631 3583 635 3587 1 cinnot
rlabel pdcontact 602 3584 606 3594 1 cinnot
rlabel ndcontact 602 3564 606 3569 1 cinnot
rlabel polycontact 1131 3762 1135 3766 1 p1
rlabel metal1 809 3539 820 3543 1 s0
rlabel ndcontact 805 3531 809 3536 1 s0
rlabel pdcontact 805 3551 809 3561 1 s0
rlabel polycontact 789 3539 793 3543 1 s0n
rlabel pdcontact 756 3548 760 3568 1 s0n
rlabel ndcontact 746 3523 752 3528 1 s0n
rlabel pdiffusion 746 3548 752 3568 1 orpms0
rlabel polycontact 739 3537 743 3541 1 or2s0
rlabel polycontact 749 3537 753 3541 1 or1s0
rlabel pdcontact 698 3525 702 3535 1 or1s0
rlabel ndcontact 698 3505 702 3510 1 or1s0
rlabel ndcontact 696 3571 700 3576 1 or2s0
rlabel pdcontact 696 3591 700 3601 1 or2s0
rlabel polycontact 680 3579 684 3583 1 and1ns0
rlabel pdcontact 639 3594 643 3604 1 and1ns0
rlabel ndcontact 648 3565 652 3575 1 and1ns0
rlabel ndiffusion 638 3565 644 3575 1 and1nms0
rlabel ndiffusion 640 3499 646 3509 1 and2nms0
rlabel polycontact 682 3513 686 3517 1 and2ns0
rlabel ndcontact 650 3499 654 3509 1 and2ns0
rlabel pdcontact 641 3528 645 3538 1 and2ns0
rlabel ndcontact 602 3508 606 3513 1 p0not
rlabel pdcontact 602 3528 606 3538 1 p0not
rlabel polycontact 633 3517 637 3521 1 p0not
rlabel polycontact 647 3583 651 3587 1 p0
rlabel polycontact 586 3516 590 3520 1 p0
rlabel polycontact 1155 3140 1159 3144 1 or1c2
rlabel metal1 1117 3132 1121 3144 1 or1c2
rlabel ndcontact 1106 3124 1110 3129 1 or1c2
rlabel pdcontact 1106 3144 1110 3154 1 or1c2
rlabel polycontact 1090 3132 1094 3136 1 or1c2n
rlabel metal1 1062 3124 1074 3128 1 or1c2n
rlabel ndcontact 1047 3116 1053 3121 1 or1c2n
rlabel pdcontact 1057 3141 1061 3161 1 or1c2n
rlabel polycontact 919 3095 923 3099 1 p0c0
rlabel polycontact 684 3082 688 3086 1 p0c0
rlabel metal1 649 3082 658 3086 1 p0c0
rlabel ndcontact 645 3074 649 3079 1 p0c0
rlabel pdcontact 645 3094 649 3104 1 p0c0
rlabel polycontact 629 3082 633 3086 1 p0c0n
rlabel metal1 603 3078 613 3082 1 p0c0n
rlabel ndcontact 597 3068 601 3078 1 p0c0n
rlabel pdcontact 588 3097 592 3107 1 p0c0n
rlabel ndiffusion 587 3068 593 3078 1 andnmc1
rlabel ndiffusion 921 3186 927 3196 1 and2nmc2
rlabel ndiffusion 926 3077 932 3087 1 and1nmc2
rlabel metal1 944 3087 952 3091 1 p1p0c0n
rlabel pdcontact 927 3106 931 3116 1 p1p0c0n
rlabel ndcontact 936 3077 940 3087 1 p1p0c0n
rlabel polycontact 968 3091 972 3095 1 p1p0c0n
rlabel metal1 988 3091 997 3095 1 p1p0c0
rlabel pdcontact 984 3103 988 3113 1 p1p0c0
rlabel ndcontact 984 3083 988 3088 1 p1p0c0
rlabel polycontact 1050 3130 1054 3134 1 p1p0c0
rlabel metal3 979 3200 991 3204 1 p1g0
rlabel ndcontact 931 3186 935 3196 1 p1g0n
rlabel pdcontact 922 3215 926 3225 1 p1g0n
rlabel polycontact 914 3203 918 3208 1 g0
rlabel pdiffusion 1047 3141 1053 3161 1 or1pmc2
rlabel pdiffusion 1162 3151 1168 3171 1 or2pmc2
rlabel pdcontact 1172 3151 1176 3171 1 c2n
rlabel ndcontact 1162 3126 1168 3131 1 c2n
rlabel polycontact 1205 3142 1209 3146 1 c2n
rlabel metal1 1235 3142 1247 3146 1 c2
rlabel pdcontact 1221 3154 1225 3164 1 c2
rlabel ndcontact 1221 3134 1225 3139 1 c2
rlabel polycontact 1165 3140 1169 3144 1 g1
rlabel ndcontact 750 3076 754 3081 1 c1
rlabel pdcontact 750 3096 754 3106 1 c1
rlabel polycontact 734 3084 738 3088 1 c1n
rlabel ndcontact 691 3068 697 3073 1 c1n
rlabel pdcontact 701 3093 705 3113 1 c1n
rlabel pdiffusion 691 3093 697 3113 1 orpmc1
rlabel polycontact 694 3082 698 3086 1 g0
rlabel polycontact 580 3086 584 3090 1 p0
rlabel metal3 512 3141 530 3147 1 c0
rlabel metal1 1058 2834 1075 2838 1 g1
rlabel ndcontact 1051 2826 1055 2831 1 g1
rlabel pdcontact 1051 2846 1055 2856 1 g1
rlabel polycontact 1035 2834 1039 2838 1 g1n
rlabel ndiffusion 993 2820 999 2830 1 and1nmg1
rlabel ndcontact 1003 2820 1007 2830 1 g1n
rlabel pdcontact 994 2849 998 2859 1 g1n
rlabel polycontact 1002 2838 1006 2842 1 b1
rlabel polycontact 986 2837 990 2842 1 a1
rlabel metal1 670 2813 683 2818 1 g0
rlabel ndcontact 664 2806 668 2811 1 g0
rlabel pdcontact 664 2826 668 2836 1 g0
rlabel ndiffusion 606 2800 612 2810 1 and1nmg0
rlabel ndcontact 616 2800 620 2810 1 g0n
rlabel pdcontact 607 2829 611 2839 1 g0n
rlabel polycontact 648 2814 652 2818 1 g0n
rlabel polycontact 599 2817 603 2822 1 a0
rlabel ndcontact 646 2806 650 2811 1 gnd
rlabel ndcontact 598 2800 602 2810 1 gnd
rlabel ndcontact 985 2820 989 2830 1 gnd
rlabel ndcontact 1033 2826 1037 2831 1 gnd
rlabel metal1 1027 2817 1061 2820 1 gnd
rlabel metal1 979 2813 1013 2816 1 gnd
rlabel metal1 640 2797 674 2800 1 gnd
rlabel metal1 592 2793 626 2796 1 gnd
rlabel metal1 640 2842 674 2846 1 vdd
rlabel metal1 592 2844 626 2848 1 vdd
rlabel metal1 979 2864 1013 2868 1 vdd
rlabel metal1 1027 2862 1061 2866 1 vdd
rlabel pdcontact 1033 2846 1037 2856 1 vdd
rlabel pdcontact 1003 2849 1007 2859 1 vdd
rlabel pdcontact 985 2849 989 2859 1 vdd
rlabel pdcontact 646 2826 650 2836 1 vdd
rlabel pdcontact 616 2829 620 2839 1 vdd
rlabel pdcontact 598 2829 602 2839 1 vdd
rlabel pdcontact 1154 3151 1158 3171 1 vdd
rlabel pdcontact 1039 3141 1043 3161 1 vdd
rlabel pdcontact 683 3093 687 3113 1 vdd
rlabel pdcontact 732 3096 736 3106 1 vdd
rlabel pdcontact 627 3094 631 3104 1 vdd
rlabel pdcontact 597 3097 601 3107 1 vdd
rlabel pdcontact 579 3097 583 3107 1 vdd
rlabel pdcontact 961 3212 965 3222 1 vdd
rlabel pdcontact 931 3215 935 3225 1 vdd
rlabel pdcontact 913 3215 917 3225 1 vdd
rlabel pdcontact 936 3106 940 3116 1 vdd
rlabel pdcontact 918 3106 922 3116 1 vdd
rlabel pdcontact 966 3103 970 3113 1 vdd
rlabel pdcontact 1088 3144 1092 3154 1 vdd
rlabel pdcontact 1203 3154 1207 3164 1 vdd
rlabel ndcontact 1203 3134 1207 3139 1 gnd
rlabel ndcontact 1172 3126 1176 3131 1 gnd
rlabel ndcontact 1154 3126 1158 3131 1 gnd
rlabel ndcontact 1088 3124 1092 3129 1 gnd
rlabel ndcontact 1057 3116 1061 3121 1 gnd
rlabel ndcontact 1039 3116 1043 3121 1 gnd
rlabel ndcontact 966 3083 970 3088 1 gnd
rlabel ndcontact 961 3192 965 3197 1 gnd
rlabel ndcontact 913 3186 917 3196 1 gnd
rlabel ndcontact 918 3077 922 3087 1 gnd
rlabel ndcontact 732 3076 736 3081 1 gnd
rlabel ndcontact 701 3068 705 3073 1 gnd
rlabel ndcontact 683 3068 687 3073 1 gnd
rlabel ndcontact 627 3074 631 3079 1 gnd
rlabel ndcontact 579 3068 583 3078 1 gnd
rlabel metal1 573 3061 607 3064 1 gnd
rlabel metal1 621 3065 655 3068 1 gnd
rlabel metal1 677 3059 711 3062 1 gnd
rlabel metal1 726 3067 760 3070 1 gnd
rlabel metal1 955 3183 989 3186 1 gnd
rlabel metal1 907 3179 941 3182 1 gnd
rlabel metal1 912 3070 946 3073 1 gnd
rlabel metal1 960 3074 994 3077 1 gnd
rlabel metal1 1033 3107 1067 3110 1 gnd
rlabel metal1 1082 3115 1116 3118 1 gnd
rlabel metal1 1148 3117 1182 3120 1 gnd
rlabel metal1 1197 3125 1231 3128 1 gnd
rlabel metal1 1197 3170 1231 3174 1 vdd
rlabel metal1 1148 3179 1182 3183 1 vdd
rlabel metal1 1082 3160 1116 3164 1 vdd
rlabel metal1 1033 3169 1067 3173 1 vdd
rlabel metal1 960 3119 994 3123 1 vdd
rlabel metal1 912 3121 946 3125 1 vdd
rlabel metal1 955 3228 989 3232 1 vdd
rlabel metal1 907 3230 941 3234 1 vdd
rlabel metal1 726 3112 760 3116 1 vdd
rlabel metal1 677 3121 711 3125 1 vdd
rlabel metal1 621 3110 655 3114 1 vdd
rlabel metal1 573 3112 607 3116 1 vdd
rlabel metal1 1123 3846 1157 3850 1 vdd
rlabel pdcontact 1129 3830 1133 3840 1 vdd
rlabel metal1 1169 3855 1203 3859 5 vdd
rlabel pdcontact 1175 3840 1179 3850 1 vdd
rlabel pdcontact 1193 3840 1197 3850 1 vdd
rlabel metal1 1217 3853 1251 3857 5 vdd
rlabel pdcontact 1223 3837 1227 3847 1 vdd
rlabel metal1 1123 3790 1157 3794 1 vdd
rlabel pdcontact 1129 3774 1133 3784 1 vdd
rlabel metal1 1171 3789 1205 3793 1 vdd
rlabel pdcontact 1177 3774 1181 3784 1 vdd
rlabel pdcontact 1195 3774 1199 3784 1 vdd
rlabel metal1 1219 3787 1253 3791 1 vdd
rlabel pdcontact 1225 3771 1229 3781 1 vdd
rlabel metal1 1277 3822 1311 3826 1 vdd
rlabel pdcontact 1283 3794 1287 3814 1 vdd
rlabel metal1 1326 3813 1360 3817 1 vdd
rlabel pdcontact 1332 3797 1336 3807 1 vdd
rlabel metal1 1277 3760 1311 3763 1 gnd
rlabel ndcontact 1283 3769 1287 3774 1 gnd
rlabel ndcontact 1301 3769 1305 3774 1 gnd
rlabel ndcontact 1332 3777 1336 3782 1 gnd
rlabel metal1 1326 3768 1360 3771 1 gnd
rlabel metal1 1219 3742 1253 3745 1 gnd
rlabel ndcontact 1177 3745 1181 3755 1 gnd
rlabel ndcontact 1225 3751 1229 3756 1 gnd
rlabel ndcontact 1129 3754 1133 3759 1 gnd
rlabel metal1 1123 3745 1157 3748 1 gnd
rlabel metal1 1123 3801 1157 3804 1 gnd
rlabel metal1 1169 3804 1203 3807 1 gnd
rlabel ndcontact 1129 3810 1133 3815 1 gnd
rlabel ndcontact 1175 3811 1179 3821 1 gnd
rlabel metal1 1171 3738 1202 3741 1 gnd
rlabel metal1 1217 3808 1251 3811 1 gnd
rlabel ndcontact 1223 3817 1227 3822 1 gnd
rlabel ndcontact 678 3571 682 3576 1 gnd
rlabel metal1 672 3562 706 3565 1 gnd
rlabel metal1 626 3492 657 3495 1 gnd
rlabel ndcontact 630 3565 634 3575 1 gnd
rlabel ndcontact 584 3564 588 3569 1 gnd
rlabel metal1 624 3558 658 3561 1 gnd
rlabel metal1 578 3555 612 3558 1 gnd
rlabel metal1 578 3499 612 3502 1 gnd
rlabel ndcontact 584 3508 588 3513 1 gnd
rlabel ndcontact 680 3505 684 3510 1 gnd
rlabel ndcontact 632 3499 636 3509 1 gnd
rlabel metal1 674 3496 708 3499 1 gnd
rlabel metal1 781 3522 815 3525 1 gnd
rlabel ndcontact 787 3531 791 3536 1 gnd
rlabel ndcontact 756 3523 760 3528 1 gnd
rlabel ndcontact 738 3523 742 3528 1 gnd
rlabel metal1 732 3514 766 3517 1 gnd
rlabel pdcontact 787 3551 791 3561 1 vdd
rlabel metal1 781 3567 815 3571 1 vdd
rlabel pdcontact 738 3548 742 3568 1 vdd
rlabel metal1 732 3576 766 3580 1 vdd
rlabel pdcontact 680 3525 684 3535 1 vdd
rlabel metal1 674 3541 708 3545 1 vdd
rlabel pdcontact 650 3528 654 3538 1 vdd
rlabel pdcontact 632 3528 636 3538 1 vdd
rlabel metal1 626 3543 660 3547 1 vdd
rlabel pdcontact 584 3528 588 3538 1 vdd
rlabel metal1 578 3544 612 3548 1 vdd
rlabel pdcontact 678 3591 682 3601 1 vdd
rlabel metal1 672 3607 706 3611 5 vdd
rlabel pdcontact 648 3594 652 3604 1 vdd
rlabel pdcontact 630 3594 634 3604 1 vdd
rlabel metal1 624 3609 658 3613 5 vdd
rlabel pdcontact 584 3584 588 3594 1 vdd
rlabel metal1 578 3600 612 3604 1 vdd
rlabel metal1 1159 2951 1170 2955 1 p1
rlabel ndcontact 1155 2943 1159 2948 1 p1
rlabel pdcontact 1155 2963 1159 2973 1 p1
rlabel polycontact 1139 2951 1143 2955 1 outnp1
rlabel ndcontact 1096 2935 1102 2940 1 outnp1
rlabel pdcontact 1106 2960 1110 2980 1 outnp1
rlabel pdiffusion 1096 2960 1102 2980 1 orpmp1
rlabel pdcontact 1046 3003 1050 3013 1 or2p1
rlabel ndcontact 1046 2983 1050 2988 1 or2p1
rlabel polycontact 1089 2949 1093 2953 1 or2p1
rlabel polycontact 1099 2949 1103 2953 1 or1p1
rlabel pdcontact 1048 2937 1052 2947 1 or1p1
rlabel ndcontact 1048 2917 1052 2922 1 or1p1
rlabel polycontact 1032 2925 1036 2929 1 and2np1
rlabel ndiffusion 990 2911 996 2921 1 and2nmp1
rlabel ndcontact 1000 2911 1004 2921 1 and2np1
rlabel pdcontact 991 2940 995 2950 1 and2np1
rlabel polycontact 999 2929 1003 2933 1 b1
rlabel polycontact 997 2995 1001 2999 1 a1
rlabel polycontact 1030 2991 1034 2995 1 and1np1
rlabel ndiffusion 988 2977 994 2987 1 and1nmp1
rlabel ndcontact 998 2977 1002 2987 1 and1np1
rlabel pdcontact 989 3006 993 3016 1 and1np1
rlabel pdcontact 952 2996 956 3006 1 b1not
rlabel ndcontact 952 2976 956 2981 1 b1not
rlabel polycontact 981 2995 985 2999 1 b1not
rlabel polycontact 983 2929 987 2933 1 a1not
rlabel pdcontact 952 2940 956 2950 1 a1not
rlabel ndcontact 952 2920 956 2925 1 a1not
rlabel polycontact 936 2928 940 2932 1 a1
rlabel polycontact 936 2984 940 2988 1 b1
rlabel pdcontact 803 2961 807 2971 1 p0
rlabel ndcontact 803 2941 807 2946 1 p0
rlabel polycontact 787 2949 791 2953 1 outnp0
rlabel ndcontact 744 2933 750 2938 1 outnp0
rlabel pdcontact 754 2958 758 2978 1 outnp0
rlabel pdiffusion 744 2958 750 2978 1 orpmp0
rlabel polycontact 747 2947 751 2951 1 or1p0
rlabel polycontact 737 2947 741 2951 1 or2p0
rlabel ndcontact 694 2981 698 2986 1 or2p0
rlabel pdcontact 694 3001 698 3011 1 or2p0
rlabel pdcontact 696 2935 700 2945 1 or1p0
rlabel ndcontact 696 2915 700 2920 1 or1p0
rlabel polycontact 680 2923 684 2927 1 and2np0
rlabel polycontact 678 2989 682 2993 1 and1np0
rlabel pdcontact 637 3004 641 3014 1 and1np0
rlabel ndiffusion 636 2975 642 2985 1 and1nmp0
rlabel ndcontact 646 2975 650 2985 1 and1np0
rlabel ndcontact 648 2909 652 2919 1 and2np0
rlabel pdcontact 639 2938 643 2948 1 and2np0
rlabel ndiffusion 638 2909 644 2919 1 and2nmp0
rlabel metal1 807 2949 818 2953 1 p0
rlabel polycontact 647 2927 651 2931 1 b0
rlabel polycontact 645 2993 649 2997 1 a0
rlabel polycontact 629 2993 633 2997 1 b0not
rlabel polycontact 631 2927 635 2931 1 a0not
rlabel ndcontact 600 2974 604 2979 1 b0not
rlabel ndcontact 600 2918 604 2923 1 a0not
rlabel polycontact 584 2926 588 2930 1 a0
rlabel polycontact 584 2982 588 2986 1 b0
rlabel ndcontact 676 2981 680 2986 1 gnd
rlabel metal1 670 2972 704 2975 1 gnd
rlabel metal1 624 2902 655 2905 1 gnd
rlabel pdcontact 600 2938 604 2948 1 anot
rlabel pdcontact 600 2994 604 3004 1 bnot
rlabel ndcontact 628 2975 632 2985 1 gnd
rlabel ndcontact 582 2974 586 2979 1 gnd
rlabel metal1 622 2968 656 2971 1 gnd
rlabel metal1 576 2965 610 2968 1 gnd
rlabel metal1 576 2909 610 2912 1 gnd
rlabel ndcontact 582 2918 586 2923 1 gnd
rlabel ndcontact 678 2915 682 2920 1 gnd
rlabel ndcontact 630 2909 634 2919 1 gnd
rlabel metal1 672 2906 706 2909 1 gnd
rlabel metal1 779 2932 813 2935 1 gnd
rlabel ndcontact 785 2941 789 2946 1 gnd
rlabel ndcontact 754 2933 758 2938 1 gnd
rlabel ndcontact 736 2933 740 2938 1 gnd
rlabel metal1 730 2924 764 2927 1 gnd
rlabel pdcontact 785 2961 789 2971 1 vdd
rlabel metal1 779 2977 813 2981 1 vdd
rlabel pdcontact 736 2958 740 2978 1 vdd
rlabel metal1 730 2986 764 2990 1 vdd
rlabel pdcontact 678 2935 682 2945 1 vdd
rlabel metal1 672 2951 706 2955 1 vdd
rlabel pdcontact 648 2938 652 2948 1 vdd
rlabel pdcontact 630 2938 634 2948 1 vdd
rlabel metal1 624 2953 658 2957 1 vdd
rlabel pdcontact 582 2938 586 2948 1 vdd
rlabel metal1 576 2954 610 2958 1 vdd
rlabel pdcontact 676 3001 680 3011 1 vdd
rlabel metal1 670 3017 704 3021 5 vdd
rlabel pdcontact 646 3004 650 3014 1 vdd
rlabel pdcontact 628 3004 632 3014 1 vdd
rlabel metal1 622 3019 656 3023 5 vdd
rlabel pdcontact 582 2994 586 3004 1 vdd
rlabel metal1 576 3010 610 3014 1 vdd
rlabel ndcontact 1028 2983 1032 2988 1 gnd
rlabel metal1 1022 2974 1056 2977 1 gnd
rlabel metal1 976 2904 1007 2907 1 gnd
rlabel ndcontact 980 2977 984 2987 1 gnd
rlabel ndcontact 934 2976 938 2981 1 gnd
rlabel metal1 974 2970 1008 2973 1 gnd
rlabel metal1 928 2967 962 2970 1 gnd
rlabel metal1 928 2911 962 2914 1 gnd
rlabel ndcontact 934 2920 938 2925 1 gnd
rlabel ndcontact 1030 2917 1034 2922 1 gnd
rlabel ndcontact 982 2911 986 2921 1 gnd
rlabel metal1 1024 2908 1058 2911 1 gnd
rlabel metal1 1131 2934 1165 2937 1 gnd
rlabel ndcontact 1137 2943 1141 2948 1 gnd
rlabel ndcontact 1106 2935 1110 2940 1 gnd
rlabel ndcontact 1088 2935 1092 2940 1 gnd
rlabel metal1 1082 2926 1116 2929 1 gnd
rlabel pdcontact 1137 2963 1141 2973 1 vdd
rlabel metal1 1131 2979 1165 2983 1 vdd
rlabel pdcontact 1088 2960 1092 2980 1 vdd
rlabel metal1 1082 2988 1116 2992 1 vdd
rlabel pdcontact 1030 2937 1034 2947 1 vdd
rlabel metal1 1024 2953 1058 2957 1 vdd
rlabel pdcontact 1000 2940 1004 2950 1 vdd
rlabel pdcontact 982 2940 986 2950 1 vdd
rlabel metal1 976 2955 1010 2959 1 vdd
rlabel pdcontact 934 2940 938 2950 1 vdd
rlabel metal1 928 2956 962 2960 1 vdd
rlabel pdcontact 1028 3003 1032 3013 1 vdd
rlabel metal1 1022 3019 1056 3023 5 vdd
rlabel pdcontact 998 3006 1002 3016 1 vdd
rlabel pdcontact 980 3006 984 3016 1 vdd
rlabel metal1 974 3021 1008 3025 5 vdd
rlabel pdcontact 934 2996 938 3006 1 vdd
rlabel metal1 928 3012 962 3016 1 vdd
rlabel metal1 2353 2962 2359 2966 1 outnp3
rlabel polycontact 2325 2968 2329 2972 1 or2p3
rlabel metal2 2298 2965 2307 2968 1 or1p3
rlabel metal1 2286 3010 2295 3014 1 or2p3
rlabel pdcontact 1554 3126 1558 3136 1 p2g1
rlabel ndcontact 1554 3106 1558 3111 1 p2g1
rlabel metal2 2292 2944 2303 2948 1 or1p3
rlabel metal2 2597 3803 2605 3807 1 or1s3
rlabel polycontact 596 3086 600 3090 1 c0
rlabel polycontact 1505 3118 1509 3122 1 g1
rlabel polycontact 1991 3231 1995 3235 1 g2
rlabel polysilicon 698 3082 700 3086 1 g0
rlabel polysilicon 1169 3140 1171 3144 1 g1
rlabel polysilicon 1503 3118 1505 3122 1 g1
rlabel polysilicon 1989 3231 1991 3235 1 g2
rlabel polysilicon 2485 3307 2487 3311 1 g3
rlabel polysilicon 2339 2968 2341 2972 1 or1p3
rlabel polysilicon 2641 3827 2643 3831 1 or1s3
rlabel polysilicon 594 3086 596 3090 1 c0
rlabel polysilicon 2124 3418 2126 3422 1 p3p2p1p0c0
rlabel polycontact 2119 3174 2123 3178 1 p3p2g1
rlabel polysilicon 2123 3174 2125 3178 1 p3p2g1
rlabel m3contact 545 2941 552 2946 1 b0
rlabel m3contact 524 2850 532 2856 1 a0
rlabel m3contact 887 2837 894 2842 1 a1
rlabel m3contact 1431 2930 1436 2936 1 a2
rlabel metal2 1566 2876 1571 2882 1 b2
rlabel m3contact 2150 3025 2155 3033 1 a3
rlabel polycontact 2222 2869 2226 2873 1 b3
rlabel m3contact 2236 2900 2241 2905 1 b3
rlabel metal1 761 3084 774 3089 1 c1
<< end >>
