magic
tech scmos
timestamp 1732058446
<< nwell >>
rect 4450 965 4484 991
rect 4496 975 4530 1000
rect 4544 972 4578 998
rect 4995 974 5029 1000
rect 5041 984 5075 1009
rect 5089 981 5123 1007
rect 5576 991 5610 1017
rect 5622 1001 5656 1026
rect 5670 998 5704 1024
rect 6134 993 6168 1019
rect 6180 1003 6214 1028
rect 6228 1000 6262 1026
rect 4450 909 4484 935
rect 4498 909 4532 934
rect 4546 906 4580 932
rect 4604 929 4638 967
rect 4653 932 4687 958
rect 4995 918 5029 944
rect 5043 918 5077 943
rect 5091 915 5125 941
rect 5149 938 5183 976
rect 5198 941 5232 967
rect 5576 935 5610 961
rect 5624 935 5658 960
rect 5672 932 5706 958
rect 5730 955 5764 993
rect 5779 958 5813 984
rect 6134 937 6168 963
rect 6182 937 6216 962
rect 6230 934 6264 960
rect 6288 957 6322 995
rect 6337 960 6371 986
<< ntransistor >>
rect 5588 977 5590 982
rect 5633 978 5635 988
rect 5643 978 5645 988
rect 5682 984 5684 989
rect 4462 951 4464 956
rect 4507 952 4509 962
rect 4517 952 4519 962
rect 4556 958 4558 963
rect 5007 960 5009 965
rect 5052 961 5054 971
rect 5062 961 5064 971
rect 5101 967 5103 972
rect 6146 979 6148 984
rect 6191 980 6193 990
rect 6201 980 6203 990
rect 6240 986 6242 991
rect 4462 895 4464 900
rect 4665 918 4667 923
rect 4615 910 4617 915
rect 4625 910 4627 915
rect 5007 904 5009 909
rect 5210 927 5212 932
rect 5160 919 5162 924
rect 5170 919 5172 924
rect 5588 921 5590 926
rect 5791 944 5793 949
rect 5741 936 5743 941
rect 5751 936 5753 941
rect 6146 923 6148 928
rect 6349 946 6351 951
rect 6299 938 6301 943
rect 6309 938 6311 943
rect 5635 912 5637 922
rect 5645 912 5647 922
rect 5684 918 5686 923
rect 6193 914 6195 924
rect 6203 914 6205 924
rect 6242 920 6244 925
rect 4509 886 4511 896
rect 4519 886 4521 896
rect 4558 892 4560 897
rect 5054 895 5056 905
rect 5064 895 5066 905
rect 5103 901 5105 906
<< ptransistor >>
rect 5633 1007 5635 1017
rect 5643 1007 5645 1017
rect 4507 981 4509 991
rect 4517 981 4519 991
rect 5052 990 5054 1000
rect 5062 990 5064 1000
rect 5588 997 5590 1007
rect 4462 971 4464 981
rect 4556 978 4558 988
rect 5007 980 5009 990
rect 5101 987 5103 997
rect 5682 1004 5684 1014
rect 6191 1009 6193 1019
rect 6201 1009 6203 1019
rect 6146 999 6148 1009
rect 6240 1006 6242 1016
rect 4615 935 4617 955
rect 4625 935 4627 955
rect 4665 938 4667 948
rect 5160 944 5162 964
rect 5170 944 5172 964
rect 5741 961 5743 981
rect 5751 961 5753 981
rect 5791 964 5793 974
rect 5210 947 5212 957
rect 4462 915 4464 925
rect 4509 915 4511 925
rect 4519 915 4521 925
rect 4558 912 4560 922
rect 5007 924 5009 934
rect 5054 924 5056 934
rect 5064 924 5066 934
rect 5103 921 5105 931
rect 5588 941 5590 951
rect 5635 941 5637 951
rect 5645 941 5647 951
rect 5684 938 5686 948
rect 6299 963 6301 983
rect 6309 963 6311 983
rect 6349 966 6351 976
rect 6146 943 6148 953
rect 6193 943 6195 953
rect 6203 943 6205 953
rect 6242 940 6244 950
<< ndiffusion >>
rect 5586 977 5588 982
rect 5590 977 5600 982
rect 5632 978 5633 988
rect 5635 978 5643 988
rect 5645 978 5646 988
rect 5680 984 5682 989
rect 5684 984 5694 989
rect 4460 951 4462 956
rect 4464 951 4474 956
rect 4506 952 4507 962
rect 4509 952 4517 962
rect 4519 952 4520 962
rect 4554 958 4556 963
rect 4558 958 4568 963
rect 5005 960 5007 965
rect 5009 960 5019 965
rect 5051 961 5052 971
rect 5054 961 5062 971
rect 5064 961 5065 971
rect 5099 967 5101 972
rect 5103 967 5113 972
rect 6144 979 6146 984
rect 6148 979 6158 984
rect 6190 980 6191 990
rect 6193 980 6201 990
rect 6203 980 6204 990
rect 6238 986 6240 991
rect 6242 986 6252 991
rect 4460 895 4462 900
rect 4464 895 4474 900
rect 4663 918 4665 923
rect 4667 918 4677 923
rect 4614 910 4615 915
rect 4617 910 4618 915
rect 4624 910 4625 915
rect 4627 910 4628 915
rect 5005 904 5007 909
rect 5009 904 5019 909
rect 5208 927 5210 932
rect 5212 927 5222 932
rect 5159 919 5160 924
rect 5162 919 5163 924
rect 5169 919 5170 924
rect 5172 919 5173 924
rect 5586 921 5588 926
rect 5590 921 5600 926
rect 5789 944 5791 949
rect 5793 944 5803 949
rect 5740 936 5741 941
rect 5743 936 5744 941
rect 5750 936 5751 941
rect 5753 936 5754 941
rect 6144 923 6146 928
rect 6148 923 6158 928
rect 6347 946 6349 951
rect 6351 946 6361 951
rect 6298 938 6299 943
rect 6301 938 6302 943
rect 6308 938 6309 943
rect 6311 938 6312 943
rect 5634 912 5635 922
rect 5637 912 5645 922
rect 5647 912 5648 922
rect 5682 918 5684 923
rect 5686 918 5696 923
rect 6192 914 6193 924
rect 6195 914 6203 924
rect 6205 914 6206 924
rect 6240 920 6242 925
rect 6244 920 6254 925
rect 4508 886 4509 896
rect 4511 886 4519 896
rect 4521 886 4522 896
rect 4556 892 4558 897
rect 4560 892 4570 897
rect 5053 895 5054 905
rect 5056 895 5064 905
rect 5066 895 5067 905
rect 5101 901 5103 906
rect 5105 901 5115 906
<< pdiffusion >>
rect 5632 1007 5633 1017
rect 5635 1007 5637 1017
rect 5641 1007 5643 1017
rect 5645 1007 5646 1017
rect 4506 981 4507 991
rect 4509 981 4511 991
rect 4515 981 4517 991
rect 4519 981 4520 991
rect 5051 990 5052 1000
rect 5054 990 5056 1000
rect 5060 990 5062 1000
rect 5064 990 5065 1000
rect 5586 997 5588 1007
rect 5590 997 5600 1007
rect 4460 971 4462 981
rect 4464 971 4474 981
rect 4554 978 4556 988
rect 4558 978 4568 988
rect 5005 980 5007 990
rect 5009 980 5019 990
rect 5099 987 5101 997
rect 5103 987 5113 997
rect 5680 1004 5682 1014
rect 5684 1004 5694 1014
rect 6190 1009 6191 1019
rect 6193 1009 6195 1019
rect 6199 1009 6201 1019
rect 6203 1009 6204 1019
rect 6144 999 6146 1009
rect 6148 999 6158 1009
rect 6238 1006 6240 1016
rect 6242 1006 6252 1016
rect 4614 935 4615 955
rect 4617 935 4625 955
rect 4627 935 4628 955
rect 4663 938 4665 948
rect 4667 938 4677 948
rect 5159 944 5160 964
rect 5162 944 5170 964
rect 5172 944 5173 964
rect 5740 961 5741 981
rect 5743 961 5751 981
rect 5753 961 5754 981
rect 5789 964 5791 974
rect 5793 964 5803 974
rect 5208 947 5210 957
rect 5212 947 5222 957
rect 4460 915 4462 925
rect 4464 915 4474 925
rect 4508 915 4509 925
rect 4511 915 4513 925
rect 4517 915 4519 925
rect 4521 915 4522 925
rect 4556 912 4558 922
rect 4560 912 4570 922
rect 5005 924 5007 934
rect 5009 924 5019 934
rect 5053 924 5054 934
rect 5056 924 5058 934
rect 5062 924 5064 934
rect 5066 924 5067 934
rect 5101 921 5103 931
rect 5105 921 5115 931
rect 5586 941 5588 951
rect 5590 941 5600 951
rect 5634 941 5635 951
rect 5637 941 5639 951
rect 5643 941 5645 951
rect 5647 941 5648 951
rect 5682 938 5684 948
rect 5686 938 5696 948
rect 6298 963 6299 983
rect 6301 963 6309 983
rect 6311 963 6312 983
rect 6347 966 6349 976
rect 6351 966 6361 976
rect 6144 943 6146 953
rect 6148 943 6158 953
rect 6192 943 6193 953
rect 6195 943 6197 953
rect 6201 943 6203 953
rect 6205 943 6206 953
rect 6240 940 6242 950
rect 6244 940 6254 950
<< ndcontact >>
rect 5582 977 5586 982
rect 5600 977 5604 982
rect 5628 978 5632 988
rect 5646 978 5650 988
rect 5676 984 5680 989
rect 5694 984 5698 989
rect 4456 951 4460 956
rect 4474 951 4478 956
rect 4502 952 4506 962
rect 4520 952 4524 962
rect 4550 958 4554 963
rect 4568 958 4572 963
rect 5001 960 5005 965
rect 5019 960 5023 965
rect 5047 961 5051 971
rect 5065 961 5069 971
rect 5095 967 5099 972
rect 5113 967 5117 972
rect 6140 979 6144 984
rect 6158 979 6162 984
rect 6186 980 6190 990
rect 6204 980 6208 990
rect 6234 986 6238 991
rect 6252 986 6256 991
rect 4456 895 4460 900
rect 4474 895 4478 900
rect 4659 918 4663 923
rect 4677 918 4681 923
rect 4610 910 4614 915
rect 4618 910 4624 915
rect 4628 910 4632 915
rect 5001 904 5005 909
rect 5019 904 5023 909
rect 5204 927 5208 932
rect 5222 927 5226 932
rect 5155 919 5159 924
rect 5163 919 5169 924
rect 5173 919 5177 924
rect 5582 921 5586 926
rect 5600 921 5604 926
rect 5785 944 5789 949
rect 5803 944 5807 949
rect 5736 936 5740 941
rect 5744 936 5750 941
rect 5754 936 5758 941
rect 6140 923 6144 928
rect 6158 923 6162 928
rect 6343 946 6347 951
rect 6361 946 6365 951
rect 6294 938 6298 943
rect 6302 938 6308 943
rect 6312 938 6316 943
rect 5630 912 5634 922
rect 5648 912 5652 922
rect 5678 918 5682 923
rect 5696 918 5700 923
rect 6188 914 6192 924
rect 6206 914 6210 924
rect 6236 920 6240 925
rect 6254 920 6258 925
rect 4504 886 4508 896
rect 4522 886 4526 896
rect 4552 892 4556 897
rect 4570 892 4574 897
rect 5049 895 5053 905
rect 5067 895 5071 905
rect 5097 901 5101 906
rect 5115 901 5119 906
<< pdcontact >>
rect 5628 1007 5632 1017
rect 5637 1007 5641 1017
rect 5646 1007 5650 1017
rect 4502 981 4506 991
rect 4511 981 4515 991
rect 4520 981 4524 991
rect 5047 990 5051 1000
rect 5056 990 5060 1000
rect 5065 990 5069 1000
rect 5582 997 5586 1007
rect 5600 997 5604 1007
rect 4456 971 4460 981
rect 4474 971 4478 981
rect 4550 978 4554 988
rect 4568 978 4572 988
rect 5001 980 5005 990
rect 5019 980 5023 990
rect 5095 987 5099 997
rect 5113 987 5117 997
rect 5676 1004 5680 1014
rect 5694 1004 5698 1014
rect 6186 1009 6190 1019
rect 6195 1009 6199 1019
rect 6204 1009 6208 1019
rect 6140 999 6144 1009
rect 6158 999 6162 1009
rect 6234 1006 6238 1016
rect 6252 1006 6256 1016
rect 4610 935 4614 955
rect 4628 935 4632 955
rect 4659 938 4663 948
rect 4677 938 4681 948
rect 5155 944 5159 964
rect 5173 944 5177 964
rect 5736 961 5740 981
rect 5754 961 5758 981
rect 5785 964 5789 974
rect 5803 964 5807 974
rect 5204 947 5208 957
rect 5222 947 5226 957
rect 4456 915 4460 925
rect 4474 915 4478 925
rect 4504 915 4508 925
rect 4513 915 4517 925
rect 4522 915 4526 925
rect 4552 912 4556 922
rect 4570 912 4574 922
rect 5001 924 5005 934
rect 5019 924 5023 934
rect 5049 924 5053 934
rect 5058 924 5062 934
rect 5067 924 5071 934
rect 5097 921 5101 931
rect 5115 921 5119 931
rect 5582 941 5586 951
rect 5600 941 5604 951
rect 5630 941 5634 951
rect 5639 941 5643 951
rect 5648 941 5652 951
rect 5678 938 5682 948
rect 5696 938 5700 948
rect 6294 963 6298 983
rect 6312 963 6316 983
rect 6343 966 6347 976
rect 6361 966 6365 976
rect 6140 943 6144 953
rect 6158 943 6162 953
rect 6188 943 6192 953
rect 6197 943 6201 953
rect 6206 943 6210 953
rect 6236 940 6240 950
rect 6254 940 6258 950
<< polysilicon >>
rect 5633 1017 5635 1020
rect 5643 1017 5645 1020
rect 6191 1019 6193 1022
rect 6201 1019 6203 1022
rect 5588 1007 5590 1010
rect 5682 1014 5684 1017
rect 5052 1000 5054 1003
rect 5062 1000 5064 1003
rect 4507 991 4509 994
rect 4517 991 4519 994
rect 4462 981 4464 984
rect 4556 988 4558 991
rect 5007 990 5009 993
rect 5101 997 5103 1000
rect 4462 956 4464 971
rect 4507 962 4509 981
rect 4517 962 4519 981
rect 4556 963 4558 978
rect 5007 965 5009 980
rect 5052 971 5054 990
rect 5062 971 5064 990
rect 5101 972 5103 987
rect 5588 982 5590 997
rect 5633 988 5635 1007
rect 5643 988 5645 1007
rect 6146 1009 6148 1012
rect 6240 1016 6242 1019
rect 5682 989 5684 1004
rect 6146 984 6148 999
rect 6191 990 6193 1009
rect 6201 990 6203 1009
rect 6240 991 6242 1006
rect 5682 981 5684 984
rect 5741 981 5743 984
rect 5751 981 5753 984
rect 5588 974 5590 977
rect 5633 975 5635 978
rect 5643 975 5645 978
rect 5101 964 5103 967
rect 5160 964 5162 967
rect 5170 964 5172 967
rect 4556 955 4558 958
rect 4615 955 4617 958
rect 4625 955 4627 958
rect 5007 957 5009 960
rect 5052 958 5054 961
rect 5062 958 5064 961
rect 4462 948 4464 951
rect 4507 949 4509 952
rect 4517 949 4519 952
rect 4665 948 4667 951
rect 6240 983 6242 986
rect 6299 983 6301 986
rect 6309 983 6311 986
rect 5791 974 5793 977
rect 6146 976 6148 979
rect 6191 977 6193 980
rect 6201 977 6203 980
rect 5210 957 5212 960
rect 5588 951 5590 954
rect 5635 951 5637 954
rect 5645 951 5647 954
rect 4462 925 4464 928
rect 4509 925 4511 928
rect 4519 925 4521 928
rect 4558 922 4560 925
rect 4462 900 4464 915
rect 4509 896 4511 915
rect 4519 896 4521 915
rect 4615 915 4617 935
rect 4625 915 4627 935
rect 4665 923 4667 938
rect 5007 934 5009 937
rect 5054 934 5056 937
rect 5064 934 5066 937
rect 5103 931 5105 934
rect 4665 915 4667 918
rect 4558 897 4560 912
rect 4615 907 4617 910
rect 4625 907 4627 910
rect 5007 909 5009 924
rect 5054 905 5056 924
rect 5064 905 5066 924
rect 5160 924 5162 944
rect 5170 924 5172 944
rect 5210 932 5212 947
rect 5684 948 5686 951
rect 5210 924 5212 927
rect 5588 926 5590 941
rect 5103 906 5105 921
rect 5635 922 5637 941
rect 5645 922 5647 941
rect 5741 941 5743 961
rect 5751 941 5753 961
rect 5791 949 5793 964
rect 6349 976 6351 979
rect 6146 953 6148 956
rect 6193 953 6195 956
rect 6203 953 6205 956
rect 5791 941 5793 944
rect 6242 950 6244 953
rect 5684 923 5686 938
rect 5741 933 5743 936
rect 5751 933 5753 936
rect 6146 928 6148 943
rect 6193 924 6195 943
rect 6203 924 6205 943
rect 6299 943 6301 963
rect 6309 943 6311 963
rect 6349 951 6351 966
rect 6349 943 6351 946
rect 6242 925 6244 940
rect 6299 935 6301 938
rect 6309 935 6311 938
rect 5160 916 5162 919
rect 5170 916 5172 919
rect 5588 918 5590 921
rect 6146 920 6148 923
rect 5684 915 5686 918
rect 6242 917 6244 920
rect 5635 909 5637 912
rect 5645 909 5647 912
rect 6193 911 6195 914
rect 6203 911 6205 914
rect 5007 901 5009 904
rect 4462 892 4464 895
rect 5103 898 5105 901
rect 5054 892 5056 895
rect 5064 892 5066 895
rect 4558 889 4560 892
rect 4509 883 4511 886
rect 4519 883 4521 886
<< polycontact >>
rect 4458 959 4462 963
rect 4503 970 4507 974
rect 4519 970 4523 974
rect 4552 966 4556 970
rect 5003 968 5007 972
rect 5048 979 5052 983
rect 5064 979 5068 983
rect 5097 975 5101 979
rect 5584 985 5588 989
rect 5629 996 5633 1000
rect 5645 996 5649 1000
rect 5678 992 5682 996
rect 6142 987 6146 991
rect 6187 998 6191 1002
rect 6203 998 6207 1002
rect 6236 994 6240 998
rect 4611 924 4615 928
rect 4458 903 4462 907
rect 4505 904 4509 908
rect 4621 924 4625 928
rect 4661 926 4665 930
rect 5156 933 5160 937
rect 4521 904 4525 908
rect 4554 900 4558 904
rect 5003 912 5007 916
rect 5050 913 5054 917
rect 5166 933 5170 937
rect 5206 935 5210 939
rect 5737 950 5741 954
rect 5584 929 5588 933
rect 5631 930 5635 934
rect 5066 913 5070 917
rect 5099 909 5103 913
rect 5747 950 5751 954
rect 5787 952 5791 956
rect 6295 952 6299 956
rect 5647 930 5651 934
rect 5680 926 5684 930
rect 6142 931 6146 935
rect 6189 932 6193 936
rect 6305 952 6309 956
rect 6345 954 6349 958
rect 6205 932 6209 936
rect 6238 928 6242 932
<< metal1 >>
rect 5622 1022 5656 1026
rect 6180 1024 6214 1028
rect 5628 1017 5632 1022
rect 5646 1017 5650 1022
rect 5670 1020 5704 1024
rect 5576 1013 5610 1017
rect 5041 1005 5075 1009
rect 5582 1007 5586 1013
rect 5676 1014 5680 1020
rect 6186 1019 6190 1024
rect 6204 1019 6208 1024
rect 6228 1022 6262 1026
rect 6134 1015 6168 1019
rect 5047 1000 5051 1005
rect 5065 1000 5069 1005
rect 5089 1003 5123 1007
rect 4496 996 4530 1000
rect 4502 991 4506 996
rect 4520 991 4524 996
rect 4544 994 4578 998
rect 4995 996 5029 1000
rect 4450 987 4484 991
rect 4456 981 4460 987
rect 4550 988 4554 994
rect 5001 990 5005 996
rect 5095 997 5099 1003
rect 5541 998 5561 1005
rect 4426 963 4429 964
rect 4474 963 4478 971
rect 4487 970 4503 974
rect 4487 963 4491 970
rect 4511 967 4515 981
rect 4958 983 4980 988
rect 4523 970 4527 974
rect 4568 970 4572 978
rect 4511 966 4524 967
rect 4537 966 4552 970
rect 4568 966 4588 970
rect 4971 972 4974 973
rect 5019 972 5023 980
rect 5032 979 5048 983
rect 5032 972 5036 979
rect 5056 976 5060 990
rect 5068 979 5072 983
rect 5113 979 5117 987
rect 5552 989 5555 990
rect 5600 989 5604 997
rect 5613 996 5629 1000
rect 5613 989 5617 996
rect 5637 993 5641 1007
rect 5649 996 5653 1000
rect 5694 996 5698 1004
rect 6140 1009 6144 1015
rect 6234 1016 6238 1022
rect 5637 992 5650 993
rect 5663 992 5678 996
rect 5694 992 5714 996
rect 5637 989 5667 992
rect 5694 989 5698 992
rect 5552 985 5584 989
rect 5600 985 5617 989
rect 5646 988 5667 989
rect 5600 982 5604 985
rect 5056 975 5069 976
rect 5082 975 5097 979
rect 5113 975 5133 979
rect 5676 978 5680 984
rect 5056 972 5086 975
rect 5113 972 5117 975
rect 4971 968 5003 972
rect 5019 968 5036 972
rect 5065 971 5086 972
rect 4511 963 4541 966
rect 4568 963 4572 966
rect 4426 959 4458 963
rect 4474 959 4491 963
rect 4520 962 4541 963
rect 4474 956 4478 959
rect 4550 952 4554 958
rect 4456 945 4460 951
rect 4502 948 4506 952
rect 4544 949 4578 952
rect 4496 945 4530 948
rect 4450 942 4484 945
rect 4450 931 4484 935
rect 4456 925 4460 931
rect 4498 930 4532 934
rect 4504 925 4508 930
rect 4522 925 4526 930
rect 4546 928 4580 932
rect 4583 928 4588 966
rect 4604 963 4638 967
rect 5019 965 5023 968
rect 4610 955 4614 963
rect 5095 961 5099 967
rect 4653 954 4687 958
rect 5001 954 5005 960
rect 5047 957 5051 961
rect 5089 958 5123 961
rect 5041 954 5075 957
rect 4659 948 4663 954
rect 4995 951 5029 954
rect 4995 940 5029 944
rect 4552 922 4556 928
rect 4583 924 4611 928
rect 4628 922 4632 935
rect 4677 931 4681 938
rect 5001 934 5005 940
rect 5043 939 5077 943
rect 5049 934 5053 939
rect 5067 934 5071 939
rect 5091 937 5125 941
rect 5128 937 5133 975
rect 5149 972 5183 976
rect 5155 964 5159 972
rect 5582 971 5586 977
rect 5628 974 5632 978
rect 5670 975 5704 978
rect 5622 971 5656 974
rect 5576 968 5610 971
rect 5198 963 5232 967
rect 5204 957 5208 963
rect 5576 957 5610 961
rect 4641 926 4661 930
rect 4677 926 4723 931
rect 4641 922 4645 926
rect 4677 923 4681 926
rect 5097 931 5101 937
rect 5128 933 5156 937
rect 5173 931 5177 944
rect 5222 940 5226 947
rect 5582 951 5586 957
rect 5624 956 5658 960
rect 5630 951 5634 956
rect 5648 951 5652 956
rect 5672 954 5706 958
rect 5709 954 5714 992
rect 5730 989 5764 993
rect 5736 981 5740 989
rect 6110 991 6113 992
rect 6158 991 6162 999
rect 6171 998 6187 1002
rect 6171 991 6175 998
rect 6195 995 6199 1009
rect 6207 998 6211 1002
rect 6252 998 6256 1006
rect 6195 994 6208 995
rect 6221 994 6236 998
rect 6252 994 6272 998
rect 6195 991 6225 994
rect 6252 991 6256 994
rect 6110 987 6142 991
rect 6158 987 6175 991
rect 6204 990 6225 991
rect 6158 984 6162 987
rect 5779 980 5813 984
rect 5785 974 5789 980
rect 6234 980 6238 986
rect 6140 973 6144 979
rect 6186 976 6190 980
rect 6228 977 6262 980
rect 6180 973 6214 976
rect 6134 970 6168 973
rect 5678 948 5682 954
rect 5709 950 5737 954
rect 5754 948 5758 961
rect 5803 957 5807 964
rect 6134 959 6168 963
rect 5767 952 5787 956
rect 5803 952 5824 957
rect 6140 953 6144 959
rect 6182 958 6216 962
rect 6188 953 6192 958
rect 6206 953 6210 958
rect 6230 956 6264 960
rect 6267 956 6272 994
rect 6288 991 6322 995
rect 6294 983 6298 991
rect 6337 982 6371 986
rect 6343 976 6347 982
rect 5767 948 5771 952
rect 5803 949 5807 952
rect 5186 935 5206 939
rect 5222 935 5239 940
rect 5186 931 5190 935
rect 5222 932 5226 935
rect 4474 907 4478 915
rect 4488 907 4505 908
rect 4442 903 4458 907
rect 4474 904 4505 907
rect 4474 903 4489 904
rect 4474 900 4478 903
rect 4513 901 4517 915
rect 4628 921 4645 922
rect 4618 918 4645 921
rect 4618 915 4624 918
rect 4525 904 4529 908
rect 4570 904 4574 912
rect 4659 912 4663 918
rect 5019 916 5023 924
rect 5033 916 5050 917
rect 4987 912 5003 916
rect 5019 913 5050 916
rect 5019 912 5034 913
rect 4513 900 4526 901
rect 4539 900 4554 904
rect 4570 900 4584 904
rect 4610 904 4614 910
rect 4628 904 4632 910
rect 4653 909 4687 912
rect 5019 909 5023 912
rect 5058 910 5062 924
rect 5173 930 5190 931
rect 5163 927 5190 930
rect 5600 933 5604 941
rect 5614 933 5631 934
rect 5568 929 5584 933
rect 5600 930 5631 933
rect 5600 929 5615 930
rect 5163 924 5169 927
rect 5070 913 5074 917
rect 5115 913 5119 921
rect 5204 921 5208 927
rect 5600 926 5604 929
rect 5639 927 5643 941
rect 5754 947 5771 948
rect 5744 944 5771 947
rect 5744 941 5750 944
rect 5651 930 5655 934
rect 5696 930 5700 938
rect 5785 938 5789 944
rect 6236 950 6240 956
rect 6267 952 6295 956
rect 6312 950 6316 963
rect 6361 959 6365 966
rect 6325 954 6345 958
rect 6361 954 6384 959
rect 6325 950 6329 954
rect 6361 951 6365 954
rect 5639 926 5652 927
rect 5665 926 5680 930
rect 5696 926 5710 930
rect 5736 930 5740 936
rect 5754 930 5758 936
rect 5779 935 5813 938
rect 6158 935 6162 943
rect 6172 935 6189 936
rect 6126 931 6142 935
rect 6158 932 6189 935
rect 6158 931 6173 932
rect 5730 927 5764 930
rect 6158 928 6162 931
rect 5639 923 5669 926
rect 5696 923 5700 926
rect 5648 922 5669 923
rect 5058 909 5071 910
rect 5084 909 5099 913
rect 5115 909 5129 913
rect 5155 913 5159 919
rect 5173 913 5177 919
rect 5198 918 5232 921
rect 5582 915 5586 921
rect 5149 910 5183 913
rect 5576 912 5610 915
rect 6197 929 6201 943
rect 6312 949 6329 950
rect 6302 946 6329 949
rect 6302 943 6308 946
rect 6343 940 6347 946
rect 6209 932 6213 936
rect 6294 932 6298 938
rect 6312 932 6316 938
rect 6337 937 6371 940
rect 6197 928 6210 929
rect 6223 928 6238 932
rect 6288 929 6322 932
rect 6197 925 6227 928
rect 6206 924 6227 925
rect 5678 912 5682 918
rect 6140 917 6144 923
rect 6134 914 6168 917
rect 6236 914 6240 920
rect 5058 906 5088 909
rect 5115 906 5119 909
rect 5630 908 5634 912
rect 5672 909 5706 912
rect 6188 910 6192 914
rect 6230 911 6264 914
rect 5067 905 5088 906
rect 4604 901 4638 904
rect 4513 897 4543 900
rect 4570 897 4574 900
rect 5001 898 5005 904
rect 4522 896 4543 897
rect 4456 889 4460 895
rect 4450 886 4484 889
rect 4995 895 5029 898
rect 5624 905 5655 908
rect 6182 907 6213 910
rect 5097 895 5101 901
rect 4552 886 4556 892
rect 5049 891 5053 895
rect 5091 892 5125 895
rect 5043 888 5074 891
rect 4504 882 4508 886
rect 4546 883 4580 886
rect 4498 879 4529 882
<< m2contact >>
rect 5561 998 5568 1005
rect 4421 959 4426 964
rect 4980 983 4987 988
rect 4527 969 4532 974
rect 4966 968 4971 973
rect 5072 978 5077 983
rect 5547 985 5552 990
rect 5653 995 5658 1000
rect 4723 926 4732 931
rect 6105 987 6110 992
rect 6211 997 6216 1002
rect 5824 952 5829 957
rect 5239 935 5246 940
rect 4435 903 4442 908
rect 4529 903 4534 908
rect 4980 912 4987 917
rect 4584 900 4589 905
rect 5561 929 5568 934
rect 5074 912 5079 917
rect 5655 929 5660 934
rect 6384 954 6390 959
rect 5710 926 5715 931
rect 6119 931 6126 936
rect 5129 909 5134 914
rect 6213 931 6218 936
<< metal2 >>
rect 5561 1030 5662 1034
rect 4980 1013 5081 1017
rect 4435 1004 4536 1008
rect 4435 976 4442 1004
rect 4405 971 4442 976
rect 4421 878 4426 959
rect 4435 908 4442 971
rect 4532 969 4536 1004
rect 4980 988 4987 1013
rect 4723 931 4732 943
rect 4619 924 4625 928
rect 4584 921 4622 924
rect 4529 878 4534 903
rect 4584 905 4589 921
rect 4966 901 4971 968
rect 4980 917 4987 983
rect 5077 978 5081 1013
rect 5561 1005 5568 1030
rect 5239 940 5246 982
rect 5164 933 5170 937
rect 5129 930 5167 933
rect 4966 887 4971 891
rect 5074 887 5079 912
rect 5129 914 5134 930
rect 5547 904 5552 985
rect 5561 934 5568 998
rect 5658 995 5662 1030
rect 6119 1032 6220 1036
rect 6119 1025 6126 1032
rect 6102 987 6105 992
rect 5824 957 5829 986
rect 5744 950 5747 954
rect 5710 947 5747 950
rect 5655 904 5660 929
rect 5710 931 5715 947
rect 5547 898 5599 904
rect 5605 898 5660 904
rect 6102 906 6110 987
rect 6119 936 6126 1020
rect 6216 997 6220 1032
rect 6384 959 6390 994
rect 6302 952 6305 956
rect 6268 949 6305 952
rect 6213 906 6218 931
rect 6254 932 6258 940
rect 6268 932 6273 949
rect 6254 928 6273 932
rect 6254 925 6258 928
rect 6102 901 6218 906
rect 4966 881 5079 887
rect 4427 872 4534 878
<< m3contact >>
rect 4966 891 4971 901
rect 6119 1020 6126 1025
rect 5599 898 5605 904
rect 4421 872 4427 878
<< metal3 >>
rect 6115 1020 6119 1025
rect 4958 891 4966 901
rect 5599 885 5605 898
rect 4405 872 4421 878
<< labels >>
rlabel polycontact 4458 959 4462 963 1 c0
rlabel polycontact 4521 904 4525 908 1 c0
rlabel polycontact 4503 970 4507 974 1 cinnot
rlabel pdcontact 4474 971 4478 981 1 cinnot
rlabel ndcontact 4474 951 4478 956 1 cinnot
rlabel metal1 4681 926 4692 930 1 s0
rlabel ndcontact 4677 918 4681 923 1 s0
rlabel pdcontact 4677 938 4681 948 1 s0
rlabel polycontact 4661 926 4665 930 1 s0n
rlabel pdcontact 4628 935 4632 955 1 s0n
rlabel ndcontact 4618 910 4624 915 1 s0n
rlabel pdiffusion 4618 935 4624 955 1 orpms0
rlabel polycontact 4611 924 4615 928 1 or2s0
rlabel polycontact 4621 924 4625 928 1 or1s0
rlabel pdcontact 4570 912 4574 922 1 or1s0
rlabel ndcontact 4570 892 4574 897 1 or1s0
rlabel ndcontact 4568 958 4572 963 1 or2s0
rlabel pdcontact 4568 978 4572 988 1 or2s0
rlabel polycontact 4552 966 4556 970 1 and1ns0
rlabel pdcontact 4511 981 4515 991 1 and1ns0
rlabel ndcontact 4520 952 4524 962 1 and1ns0
rlabel ndiffusion 4510 952 4516 962 1 and1nms0
rlabel ndiffusion 4512 886 4518 896 1 and2nms0
rlabel polycontact 4554 900 4558 904 1 and2ns0
rlabel ndcontact 4522 886 4526 896 1 and2ns0
rlabel pdcontact 4513 915 4517 925 1 and2ns0
rlabel ndcontact 4474 895 4478 900 1 p0not
rlabel pdcontact 4474 915 4478 925 1 p0not
rlabel polycontact 4505 904 4509 908 1 p0not
rlabel polycontact 4519 970 4523 974 1 p0
rlabel polycontact 4458 903 4462 907 1 p0
rlabel ndcontact 4550 958 4554 963 1 gnd
rlabel metal1 4544 949 4578 952 1 gnd
rlabel metal1 4498 879 4529 882 1 gnd
rlabel ndcontact 4502 952 4506 962 1 gnd
rlabel ndcontact 4456 951 4460 956 1 gnd
rlabel metal1 4496 945 4530 948 1 gnd
rlabel metal1 4450 942 4484 945 1 gnd
rlabel metal1 4450 886 4484 889 1 gnd
rlabel ndcontact 4456 895 4460 900 1 gnd
rlabel ndcontact 4552 892 4556 897 1 gnd
rlabel ndcontact 4504 886 4508 896 1 gnd
rlabel metal1 4546 883 4580 886 1 gnd
rlabel metal1 4653 909 4687 912 1 gnd
rlabel ndcontact 4659 918 4663 923 1 gnd
rlabel ndcontact 4628 910 4632 915 1 gnd
rlabel ndcontact 4610 910 4614 915 1 gnd
rlabel metal1 4604 901 4638 904 1 gnd
rlabel pdcontact 4659 938 4663 948 1 vdd
rlabel metal1 4653 954 4687 958 1 vdd
rlabel pdcontact 4610 935 4614 955 1 vdd
rlabel metal1 4604 963 4638 967 1 vdd
rlabel pdcontact 4552 912 4556 922 1 vdd
rlabel metal1 4546 928 4580 932 1 vdd
rlabel pdcontact 4522 915 4526 925 1 vdd
rlabel pdcontact 4504 915 4508 925 1 vdd
rlabel metal1 4498 930 4532 934 1 vdd
rlabel pdcontact 4456 915 4460 925 1 vdd
rlabel metal1 4450 931 4484 935 1 vdd
rlabel pdcontact 4550 978 4554 988 1 vdd
rlabel metal1 4544 994 4578 998 5 vdd
rlabel pdcontact 4520 981 4524 991 1 vdd
rlabel pdcontact 4502 981 4506 991 1 vdd
rlabel metal1 4496 996 4530 1000 5 vdd
rlabel pdcontact 4456 971 4460 981 1 vdd
rlabel metal1 4450 987 4484 991 1 vdd
rlabel polycontact 5064 979 5068 983 1 p1
rlabel metal1 5226 935 5237 939 1 s1
rlabel ndcontact 5222 927 5226 932 1 s1
rlabel pdcontact 5222 947 5226 957 1 s1
rlabel polycontact 5206 935 5210 939 1 s1n
rlabel ndcontact 5163 919 5169 924 1 s1n
rlabel pdcontact 5173 944 5177 964 1 s1n
rlabel pdiffusion 5163 944 5169 964 1 orpms1
rlabel pdcontact 5113 987 5117 997 1 or2s1
rlabel ndcontact 5113 967 5117 972 1 or2s1
rlabel polycontact 5166 933 5170 937 1 or1s1
rlabel polycontact 5156 933 5160 937 1 or2s1
rlabel ndcontact 5115 901 5119 906 1 or1s1
rlabel pdcontact 5115 921 5119 931 1 or1s1
rlabel ndiffusion 5057 895 5063 905 1 and2nms1
rlabel ndiffusion 5055 961 5061 971 1 and1nms1
rlabel polycontact 5097 975 5101 979 1 and1ns1
rlabel polycontact 5099 909 5103 913 1 and2ns1
rlabel ndcontact 5067 895 5071 905 1 and2ns1
rlabel ndcontact 5065 961 5069 971 1 and1ns1
rlabel pdcontact 5056 990 5060 1000 1 and1ns1
rlabel pdcontact 5058 924 5062 934 1 and2ns1
rlabel polycontact 5066 913 5070 917 1 c1
rlabel polycontact 5050 913 5054 917 1 p1not
rlabel pdcontact 5019 924 5023 934 1 p1not
rlabel ndcontact 5019 904 5023 909 1 p1not
rlabel polycontact 5048 979 5052 983 1 c1not
rlabel pdcontact 5019 980 5023 990 1 c1not
rlabel ndcontact 5019 960 5023 965 1 c1not
rlabel polycontact 5003 968 5007 972 1 c1
rlabel polycontact 5003 912 5007 916 1 p1
rlabel metal1 4995 996 5029 1000 1 vdd
rlabel pdcontact 5001 980 5005 990 1 vdd
rlabel metal1 5041 1005 5075 1009 5 vdd
rlabel pdcontact 5047 990 5051 1000 1 vdd
rlabel pdcontact 5065 990 5069 1000 1 vdd
rlabel metal1 5089 1003 5123 1007 5 vdd
rlabel pdcontact 5095 987 5099 997 1 vdd
rlabel metal1 4995 940 5029 944 1 vdd
rlabel pdcontact 5001 924 5005 934 1 vdd
rlabel metal1 5043 939 5077 943 1 vdd
rlabel pdcontact 5049 924 5053 934 1 vdd
rlabel pdcontact 5067 924 5071 934 1 vdd
rlabel metal1 5091 937 5125 941 1 vdd
rlabel pdcontact 5097 921 5101 931 1 vdd
rlabel metal1 5149 972 5183 976 1 vdd
rlabel pdcontact 5155 944 5159 964 1 vdd
rlabel metal1 5198 963 5232 967 1 vdd
rlabel pdcontact 5204 947 5208 957 1 vdd
rlabel metal1 5149 910 5183 913 1 gnd
rlabel ndcontact 5155 919 5159 924 1 gnd
rlabel ndcontact 5173 919 5177 924 1 gnd
rlabel ndcontact 5204 927 5208 932 1 gnd
rlabel metal1 5198 918 5232 921 1 gnd
rlabel metal1 5091 892 5125 895 1 gnd
rlabel ndcontact 5049 895 5053 905 1 gnd
rlabel ndcontact 5097 901 5101 906 1 gnd
rlabel ndcontact 5001 904 5005 909 1 gnd
rlabel metal1 4995 895 5029 898 1 gnd
rlabel metal1 4995 951 5029 954 1 gnd
rlabel metal1 5041 954 5075 957 1 gnd
rlabel ndcontact 5001 960 5005 965 1 gnd
rlabel ndcontact 5047 961 5051 971 1 gnd
rlabel metal1 5043 888 5074 891 1 gnd
rlabel metal1 5089 958 5123 961 1 gnd
rlabel ndcontact 5095 967 5099 972 1 gnd
rlabel metal1 5807 952 5818 956 1 s2
rlabel pdcontact 5803 964 5807 974 1 s2
rlabel ndcontact 5803 944 5807 949 1 s2
rlabel polycontact 5787 952 5791 956 1 s2n
rlabel ndcontact 5744 936 5750 941 1 s2n
rlabel pdcontact 5754 961 5758 981 1 s2n
rlabel pdiffusion 5744 961 5750 981 1 orpms2
rlabel polycontact 5747 950 5751 954 1 or1s2
rlabel pdcontact 5696 938 5700 948 1 or1s2
rlabel ndcontact 5696 918 5700 923 1 or1s2
rlabel polycontact 5737 950 5741 954 1 or2s2
rlabel ndcontact 5694 984 5698 989 1 or2s2
rlabel pdcontact 5694 1004 5698 1014 1 or2s2
rlabel polycontact 5680 926 5684 930 1 and2ns2
rlabel ndiffusion 5638 912 5644 922 1 and2nms2
rlabel ndcontact 5648 912 5652 922 1 and2ns2
rlabel pdcontact 5639 941 5643 951 1 and2ns2
rlabel polycontact 5678 992 5682 996 1 and1ns2
rlabel ndcontact 5646 978 5650 988 1 and1ns2
rlabel ndiffusion 5636 978 5642 988 1 and1nms2
rlabel pdcontact 5637 1007 5641 1017 1 and1ns2
rlabel polycontact 5629 996 5633 1000 1 p2not
rlabel pdcontact 5600 997 5604 1007 1 p2not
rlabel ndcontact 5600 977 5604 982 1 p2not
rlabel polycontact 5645 996 5649 1000 1 c2
rlabel polycontact 5584 985 5588 989 1 p2
rlabel polycontact 5647 930 5651 934 1 p2
rlabel polycontact 5631 930 5635 934 1 c2not
rlabel pdcontact 5600 941 5604 951 1 c2not
rlabel ndcontact 5600 921 5604 926 1 c2not
rlabel polycontact 5584 929 5588 933 1 c2
rlabel ndcontact 5676 984 5680 989 1 gnd
rlabel metal1 5670 975 5704 978 1 gnd
rlabel metal1 5624 905 5655 908 1 gnd
rlabel ndcontact 5628 978 5632 988 1 gnd
rlabel ndcontact 5582 977 5586 982 1 gnd
rlabel metal1 5622 971 5656 974 1 gnd
rlabel metal1 5576 968 5610 971 1 gnd
rlabel metal1 5576 912 5610 915 1 gnd
rlabel ndcontact 5582 921 5586 926 1 gnd
rlabel ndcontact 5678 918 5682 923 1 gnd
rlabel ndcontact 5630 912 5634 922 1 gnd
rlabel metal1 5672 909 5706 912 1 gnd
rlabel metal1 5779 935 5813 938 1 gnd
rlabel ndcontact 5785 944 5789 949 1 gnd
rlabel ndcontact 5754 936 5758 941 1 gnd
rlabel ndcontact 5736 936 5740 941 1 gnd
rlabel metal1 5730 927 5764 930 1 gnd
rlabel pdcontact 5785 964 5789 974 1 vdd
rlabel metal1 5779 980 5813 984 1 vdd
rlabel pdcontact 5736 961 5740 981 1 vdd
rlabel metal1 5730 989 5764 993 1 vdd
rlabel pdcontact 5678 938 5682 948 1 vdd
rlabel metal1 5672 954 5706 958 1 vdd
rlabel pdcontact 5648 941 5652 951 1 vdd
rlabel pdcontact 5630 941 5634 951 1 vdd
rlabel metal1 5624 956 5658 960 1 vdd
rlabel pdcontact 5582 941 5586 951 1 vdd
rlabel metal1 5576 957 5610 961 1 vdd
rlabel pdcontact 5676 1004 5680 1014 1 vdd
rlabel metal1 5670 1020 5704 1024 5 vdd
rlabel pdcontact 5646 1007 5650 1017 1 vdd
rlabel pdcontact 5628 1007 5632 1017 1 vdd
rlabel metal1 5622 1022 5656 1026 5 vdd
rlabel pdcontact 5582 997 5586 1007 1 vdd
rlabel metal1 5576 1013 5610 1017 1 vdd
rlabel space 6305 949 6309 956 1 or1s3
rlabel metal1 6365 954 6376 958 1 s3
rlabel ndcontact 6361 946 6365 951 1 s3
rlabel pdcontact 6361 966 6365 976 1 s3
rlabel pdiffusion 6302 963 6308 983 1 orpms3
rlabel polycontact 6345 954 6349 958 1 s3n
rlabel ndcontact 6302 938 6308 943 1 s3n
rlabel pdcontact 6312 963 6316 983 1 s3n
rlabel pdcontact 6254 940 6258 950 1 or1s3
rlabel ndcontact 6254 920 6258 925 1 or1s3
rlabel polycontact 6295 952 6299 956 1 or2s3
rlabel ndcontact 6252 986 6256 991 1 or2s3
rlabel pdcontact 6252 1006 6256 1016 1 or2s3
rlabel ndiffusion 6194 980 6200 990 1 and1nms3
rlabel ndiffusion 6196 914 6202 924 1 and2nms3
rlabel polycontact 6238 928 6242 932 1 and2ns3
rlabel ndcontact 6206 914 6210 924 1 and2ns3
rlabel pdcontact 6197 943 6201 953 1 and2ns3
rlabel polycontact 6236 994 6240 998 1 and1ns3
rlabel ndcontact 6204 980 6208 990 1 and1ns3
rlabel pdcontact 6195 1009 6199 1019 1 and1ns3
rlabel polycontact 6187 998 6191 1002 1 p3not
rlabel pdcontact 6158 999 6162 1009 1 p3not
rlabel ndcontact 6158 979 6162 984 1 p3not
rlabel polycontact 6189 932 6193 936 1 c3not
rlabel pdcontact 6158 943 6162 953 1 c3not
rlabel ndcontact 6158 923 6162 928 1 c3not
rlabel polycontact 6203 998 6207 1002 1 c3
rlabel polycontact 6142 931 6146 935 1 c3
rlabel polycontact 6205 932 6209 936 1 p3
rlabel polycontact 6142 987 6146 991 1 p3
rlabel ndcontact 6234 986 6238 991 1 gnd
rlabel metal1 6228 977 6262 980 1 gnd
rlabel metal1 6182 907 6213 910 1 gnd
rlabel ndcontact 6186 980 6190 990 1 gnd
rlabel ndcontact 6140 979 6144 984 1 gnd
rlabel metal1 6180 973 6214 976 1 gnd
rlabel metal1 6134 970 6168 973 1 gnd
rlabel metal1 6134 914 6168 917 1 gnd
rlabel ndcontact 6140 923 6144 928 1 gnd
rlabel ndcontact 6236 920 6240 925 1 gnd
rlabel ndcontact 6188 914 6192 924 1 gnd
rlabel metal1 6230 911 6264 914 1 gnd
rlabel metal1 6337 937 6371 940 1 gnd
rlabel ndcontact 6343 946 6347 951 1 gnd
rlabel ndcontact 6312 938 6316 943 1 gnd
rlabel ndcontact 6294 938 6298 943 1 gnd
rlabel metal1 6288 929 6322 932 1 gnd
rlabel pdcontact 6343 966 6347 976 1 vdd
rlabel metal1 6337 982 6371 986 1 vdd
rlabel pdcontact 6294 963 6298 983 1 vdd
rlabel metal1 6288 991 6322 995 1 vdd
rlabel pdcontact 6236 940 6240 950 1 vdd
rlabel metal1 6230 956 6264 960 1 vdd
rlabel pdcontact 6206 943 6210 953 1 vdd
rlabel pdcontact 6188 943 6192 953 1 vdd
rlabel metal1 6182 958 6216 962 1 vdd
rlabel pdcontact 6140 943 6144 953 1 vdd
rlabel metal1 6134 959 6168 963 1 vdd
rlabel pdcontact 6234 1006 6238 1016 1 vdd
rlabel metal1 6228 1022 6262 1026 5 vdd
rlabel pdcontact 6204 1009 6208 1019 1 vdd
rlabel pdcontact 6186 1009 6190 1019 1 vdd
rlabel metal1 6180 1024 6214 1028 5 vdd
rlabel pdcontact 6140 999 6144 1009 1 vdd
rlabel metal1 6134 1015 6168 1019 1 vdd
rlabel metal2 6265 928 6273 932 1 or1s3
rlabel polysilicon 6309 952 6311 956 1 or1s3
<< end >>
