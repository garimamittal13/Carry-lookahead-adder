magic
tech scmos
timestamp 1732057192
<< nwell >>
rect 2288 -81 2322 -56
rect 2336 -84 2370 -58
rect 1484 -164 1518 -139
rect 2427 -140 2461 -102
rect 2476 -137 2510 -111
rect 1532 -167 1566 -141
rect 842 -211 876 -186
rect 890 -214 924 -188
rect 1616 -212 1650 -174
rect 1665 -209 1699 -183
rect 2287 -204 2321 -179
rect 2335 -207 2369 -181
rect 350 -258 384 -233
rect 398 -261 432 -235
rect 454 -262 488 -224
rect 503 -259 537 -233
rect 968 -285 1002 -247
rect 1017 -282 1051 -256
rect 1083 -275 1117 -237
rect 1132 -272 1166 -246
rect 1483 -270 1517 -245
rect 1531 -273 1565 -247
rect 1732 -251 1766 -213
rect 1781 -248 1815 -222
rect 2603 -260 2637 -222
rect 2652 -257 2686 -231
rect 2788 -251 2822 -213
rect 2837 -248 2871 -222
rect 847 -320 881 -295
rect 895 -323 929 -297
rect 1620 -314 1654 -276
rect 1669 -311 1703 -285
rect 2292 -327 2326 -302
rect 2340 -330 2374 -304
rect 1487 -367 1521 -342
rect 1535 -370 1569 -344
rect 2426 -384 2460 -346
rect 2475 -381 2509 -355
rect 2291 -455 2325 -430
rect 2339 -458 2373 -432
<< ntransistor >>
rect 2299 -104 2301 -94
rect 2309 -104 2311 -94
rect 2348 -98 2350 -93
rect 2488 -151 2490 -146
rect 2438 -159 2440 -154
rect 2448 -159 2450 -154
rect 1495 -187 1497 -177
rect 1505 -187 1507 -177
rect 1544 -181 1546 -176
rect 853 -234 855 -224
rect 863 -234 865 -224
rect 902 -228 904 -223
rect 1677 -223 1679 -218
rect 1627 -231 1629 -226
rect 1637 -231 1639 -226
rect 2298 -227 2300 -217
rect 2308 -227 2310 -217
rect 2347 -221 2349 -216
rect 361 -281 363 -271
rect 371 -281 373 -271
rect 410 -275 412 -270
rect 515 -273 517 -268
rect 465 -281 467 -276
rect 475 -281 477 -276
rect 1144 -286 1146 -281
rect 1793 -262 1795 -257
rect 1743 -270 1745 -265
rect 1753 -270 1755 -265
rect 2849 -262 2851 -257
rect 2664 -271 2666 -266
rect 2799 -270 2801 -265
rect 2809 -270 2811 -265
rect 2614 -279 2616 -274
rect 2624 -279 2626 -274
rect 1029 -296 1031 -291
rect 1094 -294 1096 -289
rect 1104 -294 1106 -289
rect 1494 -293 1496 -283
rect 1504 -293 1506 -283
rect 1543 -287 1545 -282
rect 979 -304 981 -299
rect 989 -304 991 -299
rect 1681 -325 1683 -320
rect 858 -343 860 -333
rect 868 -343 870 -333
rect 907 -337 909 -332
rect 1631 -333 1633 -328
rect 1641 -333 1643 -328
rect 2303 -350 2305 -340
rect 2313 -350 2315 -340
rect 2352 -344 2354 -339
rect 1498 -390 1500 -380
rect 1508 -390 1510 -380
rect 1547 -384 1549 -379
rect 2487 -395 2489 -390
rect 2437 -403 2439 -398
rect 2447 -403 2449 -398
rect 2302 -478 2304 -468
rect 2312 -478 2314 -468
rect 2351 -472 2353 -467
<< ptransistor >>
rect 2299 -75 2301 -65
rect 2309 -75 2311 -65
rect 2348 -78 2350 -68
rect 2438 -134 2440 -114
rect 2448 -134 2450 -114
rect 2488 -131 2490 -121
rect 1495 -158 1497 -148
rect 1505 -158 1507 -148
rect 1544 -161 1546 -151
rect 853 -205 855 -195
rect 863 -205 865 -195
rect 902 -208 904 -198
rect 1627 -206 1629 -186
rect 1637 -206 1639 -186
rect 1677 -203 1679 -193
rect 2298 -198 2300 -188
rect 2308 -198 2310 -188
rect 2347 -201 2349 -191
rect 361 -252 363 -242
rect 371 -252 373 -242
rect 410 -255 412 -245
rect 465 -256 467 -236
rect 475 -256 477 -236
rect 515 -253 517 -243
rect 1743 -245 1745 -225
rect 1753 -245 1755 -225
rect 1793 -242 1795 -232
rect 979 -279 981 -259
rect 989 -279 991 -259
rect 1029 -276 1031 -266
rect 1094 -269 1096 -249
rect 1104 -269 1106 -249
rect 1144 -266 1146 -256
rect 1494 -264 1496 -254
rect 1504 -264 1506 -254
rect 1543 -267 1545 -257
rect 2614 -254 2616 -234
rect 2624 -254 2626 -234
rect 2664 -251 2666 -241
rect 2799 -245 2801 -225
rect 2809 -245 2811 -225
rect 2849 -242 2851 -232
rect 858 -314 860 -304
rect 868 -314 870 -304
rect 907 -317 909 -307
rect 1631 -308 1633 -288
rect 1641 -308 1643 -288
rect 1681 -305 1683 -295
rect 2303 -321 2305 -311
rect 2313 -321 2315 -311
rect 2352 -324 2354 -314
rect 1498 -361 1500 -351
rect 1508 -361 1510 -351
rect 1547 -364 1549 -354
rect 2437 -378 2439 -358
rect 2447 -378 2449 -358
rect 2487 -375 2489 -365
rect 2302 -449 2304 -439
rect 2312 -449 2314 -439
rect 2351 -452 2353 -442
<< ndiffusion >>
rect 2298 -104 2299 -94
rect 2301 -104 2309 -94
rect 2311 -104 2312 -94
rect 2346 -98 2348 -93
rect 2350 -98 2360 -93
rect 2486 -151 2488 -146
rect 2490 -151 2500 -146
rect 2437 -159 2438 -154
rect 2440 -159 2441 -154
rect 2447 -159 2448 -154
rect 2450 -159 2451 -154
rect 1494 -187 1495 -177
rect 1497 -187 1505 -177
rect 1507 -187 1508 -177
rect 1542 -181 1544 -176
rect 1546 -181 1556 -176
rect 852 -234 853 -224
rect 855 -234 863 -224
rect 865 -234 866 -224
rect 900 -228 902 -223
rect 904 -228 914 -223
rect 1675 -223 1677 -218
rect 1679 -223 1689 -218
rect 1626 -231 1627 -226
rect 1629 -231 1630 -226
rect 1636 -231 1637 -226
rect 1639 -231 1640 -226
rect 2297 -227 2298 -217
rect 2300 -227 2308 -217
rect 2310 -227 2311 -217
rect 2345 -221 2347 -216
rect 2349 -221 2359 -216
rect 360 -281 361 -271
rect 363 -281 371 -271
rect 373 -281 374 -271
rect 408 -275 410 -270
rect 412 -275 422 -270
rect 513 -273 515 -268
rect 517 -273 527 -268
rect 464 -281 465 -276
rect 467 -281 468 -276
rect 474 -281 475 -276
rect 477 -281 478 -276
rect 1142 -286 1144 -281
rect 1146 -286 1156 -281
rect 1791 -262 1793 -257
rect 1795 -262 1805 -257
rect 1742 -270 1743 -265
rect 1745 -270 1746 -265
rect 1752 -270 1753 -265
rect 1755 -270 1756 -265
rect 2847 -262 2849 -257
rect 2851 -262 2861 -257
rect 2662 -271 2664 -266
rect 2666 -271 2676 -266
rect 2798 -270 2799 -265
rect 2801 -270 2802 -265
rect 2808 -270 2809 -265
rect 2811 -270 2812 -265
rect 2613 -279 2614 -274
rect 2616 -279 2617 -274
rect 2623 -279 2624 -274
rect 2626 -279 2627 -274
rect 1027 -296 1029 -291
rect 1031 -296 1041 -291
rect 1093 -294 1094 -289
rect 1096 -294 1097 -289
rect 1103 -294 1104 -289
rect 1106 -294 1107 -289
rect 1493 -293 1494 -283
rect 1496 -293 1504 -283
rect 1506 -293 1507 -283
rect 1541 -287 1543 -282
rect 1545 -287 1555 -282
rect 978 -304 979 -299
rect 981 -304 982 -299
rect 988 -304 989 -299
rect 991 -304 992 -299
rect 1679 -325 1681 -320
rect 1683 -325 1693 -320
rect 857 -343 858 -333
rect 860 -343 868 -333
rect 870 -343 871 -333
rect 905 -337 907 -332
rect 909 -337 919 -332
rect 1630 -333 1631 -328
rect 1633 -333 1634 -328
rect 1640 -333 1641 -328
rect 1643 -333 1644 -328
rect 2302 -350 2303 -340
rect 2305 -350 2313 -340
rect 2315 -350 2316 -340
rect 2350 -344 2352 -339
rect 2354 -344 2364 -339
rect 1497 -390 1498 -380
rect 1500 -390 1508 -380
rect 1510 -390 1511 -380
rect 1545 -384 1547 -379
rect 1549 -384 1559 -379
rect 2485 -395 2487 -390
rect 2489 -395 2499 -390
rect 2436 -403 2437 -398
rect 2439 -403 2440 -398
rect 2446 -403 2447 -398
rect 2449 -403 2450 -398
rect 2301 -478 2302 -468
rect 2304 -478 2312 -468
rect 2314 -478 2315 -468
rect 2349 -472 2351 -467
rect 2353 -472 2363 -467
<< pdiffusion >>
rect 2298 -75 2299 -65
rect 2301 -75 2303 -65
rect 2307 -75 2309 -65
rect 2311 -75 2312 -65
rect 2346 -78 2348 -68
rect 2350 -78 2360 -68
rect 2437 -134 2438 -114
rect 2440 -134 2448 -114
rect 2450 -134 2451 -114
rect 2486 -131 2488 -121
rect 2490 -131 2500 -121
rect 1494 -158 1495 -148
rect 1497 -158 1499 -148
rect 1503 -158 1505 -148
rect 1507 -158 1508 -148
rect 1542 -161 1544 -151
rect 1546 -161 1556 -151
rect 852 -205 853 -195
rect 855 -205 857 -195
rect 861 -205 863 -195
rect 865 -205 866 -195
rect 900 -208 902 -198
rect 904 -208 914 -198
rect 1626 -206 1627 -186
rect 1629 -206 1637 -186
rect 1639 -206 1640 -186
rect 1675 -203 1677 -193
rect 1679 -203 1689 -193
rect 2297 -198 2298 -188
rect 2300 -198 2302 -188
rect 2306 -198 2308 -188
rect 2310 -198 2311 -188
rect 2345 -201 2347 -191
rect 2349 -201 2359 -191
rect 360 -252 361 -242
rect 363 -252 365 -242
rect 369 -252 371 -242
rect 373 -252 374 -242
rect 408 -255 410 -245
rect 412 -255 422 -245
rect 464 -256 465 -236
rect 467 -256 475 -236
rect 477 -256 478 -236
rect 513 -253 515 -243
rect 517 -253 527 -243
rect 1742 -245 1743 -225
rect 1745 -245 1753 -225
rect 1755 -245 1756 -225
rect 1791 -242 1793 -232
rect 1795 -242 1805 -232
rect 978 -279 979 -259
rect 981 -279 989 -259
rect 991 -279 992 -259
rect 1027 -276 1029 -266
rect 1031 -276 1041 -266
rect 1093 -269 1094 -249
rect 1096 -269 1104 -249
rect 1106 -269 1107 -249
rect 1142 -266 1144 -256
rect 1146 -266 1156 -256
rect 1493 -264 1494 -254
rect 1496 -264 1498 -254
rect 1502 -264 1504 -254
rect 1506 -264 1507 -254
rect 1541 -267 1543 -257
rect 1545 -267 1555 -257
rect 2613 -254 2614 -234
rect 2616 -254 2624 -234
rect 2626 -254 2627 -234
rect 2662 -251 2664 -241
rect 2666 -251 2676 -241
rect 2798 -245 2799 -225
rect 2801 -245 2809 -225
rect 2811 -245 2812 -225
rect 2847 -242 2849 -232
rect 2851 -242 2861 -232
rect 857 -314 858 -304
rect 860 -314 862 -304
rect 866 -314 868 -304
rect 870 -314 871 -304
rect 905 -317 907 -307
rect 909 -317 919 -307
rect 1630 -308 1631 -288
rect 1633 -308 1641 -288
rect 1643 -308 1644 -288
rect 1679 -305 1681 -295
rect 1683 -305 1693 -295
rect 2302 -321 2303 -311
rect 2305 -321 2307 -311
rect 2311 -321 2313 -311
rect 2315 -321 2316 -311
rect 2350 -324 2352 -314
rect 2354 -324 2364 -314
rect 1497 -361 1498 -351
rect 1500 -361 1502 -351
rect 1506 -361 1508 -351
rect 1510 -361 1511 -351
rect 1545 -364 1547 -354
rect 1549 -364 1559 -354
rect 2436 -378 2437 -358
rect 2439 -378 2447 -358
rect 2449 -378 2450 -358
rect 2485 -375 2487 -365
rect 2489 -375 2499 -365
rect 2301 -449 2302 -439
rect 2304 -449 2306 -439
rect 2310 -449 2312 -439
rect 2314 -449 2315 -439
rect 2349 -452 2351 -442
rect 2353 -452 2363 -442
<< ndcontact >>
rect 2294 -104 2298 -94
rect 2312 -104 2316 -94
rect 2342 -98 2346 -93
rect 2360 -98 2364 -93
rect 2482 -151 2486 -146
rect 2500 -151 2504 -146
rect 2433 -159 2437 -154
rect 2441 -159 2447 -154
rect 2451 -159 2455 -154
rect 1490 -187 1494 -177
rect 1508 -187 1512 -177
rect 1538 -181 1542 -176
rect 1556 -181 1560 -176
rect 848 -234 852 -224
rect 866 -234 870 -224
rect 896 -228 900 -223
rect 914 -228 918 -223
rect 1671 -223 1675 -218
rect 1689 -223 1693 -218
rect 1622 -231 1626 -226
rect 1630 -231 1636 -226
rect 1640 -231 1644 -226
rect 2293 -227 2297 -217
rect 2311 -227 2315 -217
rect 2341 -221 2345 -216
rect 2359 -221 2363 -216
rect 356 -281 360 -271
rect 374 -281 378 -271
rect 404 -275 408 -270
rect 422 -275 426 -270
rect 509 -273 513 -268
rect 527 -273 531 -268
rect 460 -281 464 -276
rect 468 -281 474 -276
rect 478 -281 482 -276
rect 1138 -286 1142 -281
rect 1156 -286 1160 -281
rect 1787 -262 1791 -257
rect 1805 -262 1809 -257
rect 1738 -270 1742 -265
rect 1746 -270 1752 -265
rect 1756 -270 1760 -265
rect 2843 -262 2847 -257
rect 2861 -262 2865 -257
rect 2658 -271 2662 -266
rect 2676 -271 2680 -266
rect 2794 -270 2798 -265
rect 2802 -270 2808 -265
rect 2812 -270 2816 -265
rect 2609 -279 2613 -274
rect 2617 -279 2623 -274
rect 2627 -279 2631 -274
rect 1023 -296 1027 -291
rect 1041 -296 1045 -291
rect 1089 -294 1093 -289
rect 1097 -294 1103 -289
rect 1107 -294 1111 -289
rect 1489 -293 1493 -283
rect 1507 -293 1511 -283
rect 1537 -287 1541 -282
rect 1555 -287 1559 -282
rect 974 -304 978 -299
rect 982 -304 988 -299
rect 992 -304 996 -299
rect 1675 -325 1679 -320
rect 1693 -325 1697 -320
rect 853 -343 857 -333
rect 871 -343 875 -333
rect 901 -337 905 -332
rect 919 -337 923 -332
rect 1626 -333 1630 -328
rect 1634 -333 1640 -328
rect 1644 -333 1648 -328
rect 2298 -350 2302 -340
rect 2316 -350 2320 -340
rect 2346 -344 2350 -339
rect 2364 -344 2368 -339
rect 1493 -390 1497 -380
rect 1511 -390 1515 -380
rect 1541 -384 1545 -379
rect 1559 -384 1563 -379
rect 2481 -395 2485 -390
rect 2499 -395 2503 -390
rect 2432 -403 2436 -398
rect 2440 -403 2446 -398
rect 2450 -403 2454 -398
rect 2297 -478 2301 -468
rect 2315 -478 2319 -468
rect 2345 -472 2349 -467
rect 2363 -472 2367 -467
<< pdcontact >>
rect 2294 -75 2298 -65
rect 2303 -75 2307 -65
rect 2312 -75 2316 -65
rect 2342 -78 2346 -68
rect 2360 -78 2364 -68
rect 2433 -134 2437 -114
rect 2451 -134 2455 -114
rect 2482 -131 2486 -121
rect 2500 -131 2504 -121
rect 1490 -158 1494 -148
rect 1499 -158 1503 -148
rect 1508 -158 1512 -148
rect 1538 -161 1542 -151
rect 1556 -161 1560 -151
rect 848 -205 852 -195
rect 857 -205 861 -195
rect 866 -205 870 -195
rect 896 -208 900 -198
rect 914 -208 918 -198
rect 1622 -206 1626 -186
rect 1640 -206 1644 -186
rect 1671 -203 1675 -193
rect 1689 -203 1693 -193
rect 2293 -198 2297 -188
rect 2302 -198 2306 -188
rect 2311 -198 2315 -188
rect 2341 -201 2345 -191
rect 2359 -201 2363 -191
rect 356 -252 360 -242
rect 365 -252 369 -242
rect 374 -252 378 -242
rect 404 -255 408 -245
rect 422 -255 426 -245
rect 460 -256 464 -236
rect 478 -256 482 -236
rect 509 -253 513 -243
rect 527 -253 531 -243
rect 1738 -245 1742 -225
rect 1756 -245 1760 -225
rect 1787 -242 1791 -232
rect 1805 -242 1809 -232
rect 974 -279 978 -259
rect 992 -279 996 -259
rect 1023 -276 1027 -266
rect 1041 -276 1045 -266
rect 1089 -269 1093 -249
rect 1107 -269 1111 -249
rect 1138 -266 1142 -256
rect 1156 -266 1160 -256
rect 1489 -264 1493 -254
rect 1498 -264 1502 -254
rect 1507 -264 1511 -254
rect 1537 -267 1541 -257
rect 1555 -267 1559 -257
rect 2609 -254 2613 -234
rect 2627 -254 2631 -234
rect 2658 -251 2662 -241
rect 2676 -251 2680 -241
rect 2794 -245 2798 -225
rect 2812 -245 2816 -225
rect 2843 -242 2847 -232
rect 2861 -242 2865 -232
rect 853 -314 857 -304
rect 862 -314 866 -304
rect 871 -314 875 -304
rect 901 -317 905 -307
rect 919 -317 923 -307
rect 1626 -308 1630 -288
rect 1644 -308 1648 -288
rect 1675 -305 1679 -295
rect 1693 -305 1697 -295
rect 2298 -321 2302 -311
rect 2307 -321 2311 -311
rect 2316 -321 2320 -311
rect 2346 -324 2350 -314
rect 2364 -324 2368 -314
rect 1493 -361 1497 -351
rect 1502 -361 1506 -351
rect 1511 -361 1515 -351
rect 1541 -364 1545 -354
rect 1559 -364 1563 -354
rect 2432 -378 2436 -358
rect 2450 -378 2454 -358
rect 2481 -375 2485 -365
rect 2499 -375 2503 -365
rect 2297 -449 2301 -439
rect 2306 -449 2310 -439
rect 2315 -449 2319 -439
rect 2345 -452 2349 -442
rect 2363 -452 2367 -442
<< polysilicon >>
rect 2299 -65 2301 -62
rect 2309 -65 2311 -62
rect 2348 -68 2350 -65
rect 2299 -94 2301 -75
rect 2309 -94 2311 -75
rect 2348 -93 2350 -78
rect 2348 -101 2350 -98
rect 2299 -107 2301 -104
rect 2309 -107 2311 -104
rect 2438 -114 2440 -111
rect 2448 -114 2450 -111
rect 2488 -121 2490 -118
rect 1495 -148 1497 -145
rect 1505 -148 1507 -145
rect 1544 -151 1546 -148
rect 1495 -177 1497 -158
rect 1505 -177 1507 -158
rect 2438 -154 2440 -134
rect 2448 -154 2450 -134
rect 2488 -146 2490 -131
rect 2488 -154 2490 -151
rect 1544 -176 1546 -161
rect 2438 -162 2440 -159
rect 2448 -162 2450 -159
rect 1544 -184 1546 -181
rect 1627 -186 1629 -183
rect 1637 -186 1639 -183
rect 1495 -190 1497 -187
rect 1505 -190 1507 -187
rect 853 -195 855 -192
rect 863 -195 865 -192
rect 902 -198 904 -195
rect 853 -224 855 -205
rect 863 -224 865 -205
rect 2298 -188 2300 -185
rect 2308 -188 2310 -185
rect 1677 -193 1679 -190
rect 2347 -191 2349 -188
rect 902 -223 904 -208
rect 465 -236 467 -233
rect 475 -236 477 -233
rect 1627 -226 1629 -206
rect 1637 -226 1639 -206
rect 1677 -218 1679 -203
rect 2298 -217 2300 -198
rect 2308 -217 2310 -198
rect 2347 -216 2349 -201
rect 1677 -226 1679 -223
rect 1743 -225 1745 -222
rect 1753 -225 1755 -222
rect 902 -231 904 -228
rect 1627 -234 1629 -231
rect 1637 -234 1639 -231
rect 361 -242 363 -239
rect 371 -242 373 -239
rect 410 -245 412 -242
rect 361 -271 363 -252
rect 371 -271 373 -252
rect 410 -270 412 -255
rect 853 -237 855 -234
rect 863 -237 865 -234
rect 515 -243 517 -240
rect 2347 -224 2349 -221
rect 2799 -225 2801 -222
rect 2809 -225 2811 -222
rect 1793 -232 1795 -229
rect 2298 -230 2300 -227
rect 2308 -230 2310 -227
rect 2614 -234 2616 -231
rect 2624 -234 2626 -231
rect 1094 -249 1096 -246
rect 1104 -249 1106 -246
rect 410 -278 412 -275
rect 465 -276 467 -256
rect 475 -276 477 -256
rect 515 -268 517 -253
rect 979 -259 981 -256
rect 989 -259 991 -256
rect 515 -276 517 -273
rect 1029 -266 1031 -263
rect 1144 -256 1146 -253
rect 1494 -254 1496 -251
rect 1504 -254 1506 -251
rect 1543 -257 1545 -254
rect 361 -284 363 -281
rect 371 -284 373 -281
rect 465 -284 467 -281
rect 475 -284 477 -281
rect 979 -299 981 -279
rect 989 -299 991 -279
rect 1029 -291 1031 -276
rect 1094 -289 1096 -269
rect 1104 -289 1106 -269
rect 1144 -281 1146 -266
rect 1494 -283 1496 -264
rect 1504 -283 1506 -264
rect 1743 -265 1745 -245
rect 1753 -265 1755 -245
rect 1793 -257 1795 -242
rect 2664 -241 2666 -238
rect 2849 -232 2851 -229
rect 1793 -265 1795 -262
rect 1543 -282 1545 -267
rect 1743 -273 1745 -270
rect 1753 -273 1755 -270
rect 2614 -274 2616 -254
rect 2624 -274 2626 -254
rect 2664 -266 2666 -251
rect 2799 -265 2801 -245
rect 2809 -265 2811 -245
rect 2849 -257 2851 -242
rect 2849 -265 2851 -262
rect 2664 -274 2666 -271
rect 2799 -273 2801 -270
rect 2809 -273 2811 -270
rect 2614 -282 2616 -279
rect 2624 -282 2626 -279
rect 1144 -289 1146 -286
rect 1543 -290 1545 -287
rect 1631 -288 1633 -285
rect 1641 -288 1643 -285
rect 1029 -299 1031 -296
rect 1094 -297 1096 -294
rect 1104 -297 1106 -294
rect 1494 -296 1496 -293
rect 1504 -296 1506 -293
rect 858 -304 860 -301
rect 868 -304 870 -301
rect 907 -307 909 -304
rect 979 -307 981 -304
rect 989 -307 991 -304
rect 858 -333 860 -314
rect 868 -333 870 -314
rect 1681 -295 1683 -292
rect 907 -332 909 -317
rect 1631 -328 1633 -308
rect 1641 -328 1643 -308
rect 1681 -320 1683 -305
rect 2303 -311 2305 -308
rect 2313 -311 2315 -308
rect 2352 -314 2354 -311
rect 1681 -328 1683 -325
rect 1631 -336 1633 -333
rect 1641 -336 1643 -333
rect 907 -340 909 -337
rect 2303 -340 2305 -321
rect 2313 -340 2315 -321
rect 2352 -339 2354 -324
rect 858 -346 860 -343
rect 868 -346 870 -343
rect 1498 -351 1500 -348
rect 1508 -351 1510 -348
rect 2352 -347 2354 -344
rect 1547 -354 1549 -351
rect 2303 -353 2305 -350
rect 2313 -353 2315 -350
rect 1498 -380 1500 -361
rect 1508 -380 1510 -361
rect 2437 -358 2439 -355
rect 2447 -358 2449 -355
rect 1547 -379 1549 -364
rect 2487 -365 2489 -362
rect 1547 -387 1549 -384
rect 1498 -393 1500 -390
rect 1508 -393 1510 -390
rect 2437 -398 2439 -378
rect 2447 -398 2449 -378
rect 2487 -390 2489 -375
rect 2487 -398 2489 -395
rect 2437 -406 2439 -403
rect 2447 -406 2449 -403
rect 2302 -439 2304 -436
rect 2312 -439 2314 -436
rect 2351 -442 2353 -439
rect 2302 -468 2304 -449
rect 2312 -468 2314 -449
rect 2351 -467 2353 -452
rect 2351 -475 2353 -472
rect 2302 -481 2304 -478
rect 2312 -481 2314 -478
<< polycontact >>
rect 2295 -87 2299 -82
rect 2311 -86 2315 -82
rect 2344 -90 2348 -86
rect 2434 -145 2438 -141
rect 1491 -169 1495 -165
rect 2444 -145 2448 -141
rect 2484 -143 2488 -139
rect 1507 -169 1511 -165
rect 1540 -173 1544 -169
rect 849 -217 853 -212
rect 865 -216 869 -212
rect 898 -220 902 -216
rect 1623 -217 1627 -213
rect 1633 -217 1637 -213
rect 1673 -215 1677 -211
rect 2294 -209 2298 -205
rect 2310 -209 2314 -205
rect 2343 -213 2347 -209
rect 357 -263 361 -259
rect 373 -263 377 -259
rect 406 -267 410 -263
rect 461 -267 465 -263
rect 471 -267 475 -263
rect 511 -265 515 -261
rect 1739 -256 1743 -252
rect 975 -290 979 -286
rect 985 -290 989 -286
rect 1025 -288 1029 -284
rect 1090 -280 1094 -276
rect 1100 -280 1104 -276
rect 1140 -278 1144 -274
rect 1490 -275 1494 -271
rect 1749 -256 1753 -252
rect 1789 -254 1793 -250
rect 2610 -265 2614 -261
rect 1506 -275 1510 -271
rect 1539 -279 1543 -275
rect 2620 -265 2624 -261
rect 2660 -263 2664 -259
rect 2795 -256 2799 -252
rect 2805 -256 2809 -252
rect 2845 -254 2849 -250
rect 854 -325 858 -321
rect 870 -325 874 -321
rect 903 -329 907 -325
rect 1627 -319 1631 -315
rect 1637 -319 1641 -315
rect 1677 -317 1681 -313
rect 2299 -332 2303 -328
rect 2315 -332 2319 -328
rect 2348 -336 2352 -332
rect 1494 -372 1498 -368
rect 1510 -372 1514 -368
rect 1543 -376 1547 -372
rect 2433 -389 2437 -385
rect 2443 -389 2447 -385
rect 2483 -387 2487 -383
rect 2298 -460 2302 -456
rect 2314 -460 2318 -456
rect 2347 -464 2351 -460
<< metal1 >>
rect 2228 -56 2266 -51
rect 2288 -60 2322 -56
rect 2294 -65 2298 -60
rect 2312 -65 2316 -60
rect 2336 -62 2370 -58
rect 2342 -68 2346 -62
rect 2244 -87 2256 -82
rect 2261 -87 2295 -82
rect 1484 -143 1518 -139
rect 1490 -148 1494 -143
rect 1508 -148 1512 -143
rect 1532 -145 1566 -141
rect 1538 -151 1542 -145
rect 1455 -169 1491 -165
rect 842 -190 876 -186
rect 848 -195 852 -190
rect 866 -195 870 -190
rect 890 -192 924 -188
rect 896 -198 900 -192
rect 834 -217 849 -212
rect 857 -219 861 -205
rect 857 -220 870 -219
rect 879 -220 898 -216
rect 857 -223 882 -220
rect 866 -224 882 -223
rect 454 -228 488 -224
rect 350 -237 384 -233
rect 356 -242 360 -237
rect 374 -242 378 -237
rect 398 -239 432 -235
rect 460 -236 464 -228
rect 404 -245 408 -239
rect 344 -263 357 -259
rect 365 -266 369 -252
rect 422 -263 426 -255
rect 503 -237 537 -233
rect 896 -234 900 -228
rect 509 -243 513 -237
rect 848 -238 852 -234
rect 890 -237 924 -234
rect 842 -241 876 -238
rect 1083 -241 1117 -237
rect 968 -251 1002 -247
rect 1089 -249 1093 -241
rect 365 -267 378 -266
rect 387 -267 406 -263
rect 422 -267 461 -263
rect 365 -270 390 -267
rect 422 -270 426 -267
rect 478 -269 482 -256
rect 527 -261 531 -253
rect 974 -259 978 -251
rect 491 -265 511 -261
rect 527 -265 541 -261
rect 491 -269 495 -265
rect 527 -268 531 -265
rect 478 -270 495 -269
rect 374 -271 390 -270
rect 468 -273 495 -270
rect 404 -281 408 -275
rect 468 -276 474 -273
rect 509 -279 513 -273
rect 1017 -260 1051 -256
rect 1023 -266 1027 -260
rect 1132 -250 1166 -246
rect 1138 -256 1142 -250
rect 356 -285 360 -281
rect 398 -284 432 -281
rect 350 -288 384 -285
rect 460 -287 464 -281
rect 478 -287 482 -281
rect 503 -282 537 -279
rect 454 -290 488 -287
rect 817 -292 840 -288
rect 835 -321 840 -292
rect 992 -292 996 -279
rect 1041 -284 1045 -276
rect 1052 -280 1090 -276
rect 1052 -284 1056 -280
rect 1107 -282 1111 -269
rect 1156 -274 1160 -266
rect 1183 -274 1188 -261
rect 1120 -278 1140 -274
rect 1156 -278 1188 -274
rect 1455 -271 1461 -169
rect 1499 -172 1503 -158
rect 1556 -169 1560 -161
rect 1576 -169 1582 -138
rect 1499 -173 1512 -172
rect 1521 -173 1540 -169
rect 1556 -173 1592 -169
rect 1499 -176 1524 -173
rect 1556 -176 1560 -173
rect 1508 -177 1524 -176
rect 1538 -187 1542 -181
rect 1490 -191 1494 -187
rect 1532 -190 1566 -187
rect 1484 -194 1518 -191
rect 1588 -213 1592 -173
rect 1616 -178 1650 -174
rect 1622 -186 1626 -178
rect 1665 -187 1699 -183
rect 1671 -193 1675 -187
rect 1588 -217 1623 -213
rect 1640 -219 1644 -206
rect 1689 -211 1693 -203
rect 2244 -205 2248 -87
rect 2303 -89 2307 -75
rect 2360 -86 2364 -78
rect 2303 -90 2316 -89
rect 2325 -90 2344 -86
rect 2360 -90 2383 -86
rect 2303 -93 2328 -90
rect 2360 -93 2364 -90
rect 2312 -94 2328 -93
rect 2342 -104 2346 -98
rect 2294 -108 2298 -104
rect 2336 -107 2370 -104
rect 2288 -111 2322 -108
rect 2380 -141 2383 -90
rect 2427 -106 2461 -102
rect 2433 -114 2437 -106
rect 2476 -115 2510 -111
rect 2482 -121 2486 -115
rect 2380 -145 2434 -141
rect 2451 -147 2455 -134
rect 2500 -139 2504 -131
rect 2464 -143 2484 -139
rect 2500 -143 2564 -139
rect 2464 -147 2468 -143
rect 2500 -146 2504 -143
rect 2451 -148 2468 -147
rect 2441 -151 2468 -148
rect 2441 -154 2447 -151
rect 2482 -157 2486 -151
rect 2433 -165 2437 -159
rect 2451 -165 2455 -159
rect 2476 -160 2510 -157
rect 2427 -168 2461 -165
rect 2287 -183 2321 -179
rect 2293 -188 2297 -183
rect 2311 -188 2315 -183
rect 2335 -185 2369 -181
rect 2341 -191 2345 -185
rect 2244 -209 2294 -205
rect 1653 -215 1673 -211
rect 1689 -215 1709 -211
rect 1653 -219 1657 -215
rect 1689 -218 1693 -215
rect 1640 -220 1657 -219
rect 1630 -223 1657 -220
rect 1630 -226 1636 -223
rect 1671 -229 1675 -223
rect 1622 -237 1626 -231
rect 1640 -237 1644 -231
rect 1665 -232 1699 -229
rect 1616 -240 1650 -237
rect 1483 -249 1517 -245
rect 1489 -254 1493 -249
rect 1507 -254 1511 -249
rect 1531 -251 1565 -247
rect 1537 -257 1541 -251
rect 1706 -252 1709 -215
rect 1732 -217 1766 -213
rect 1738 -225 1742 -217
rect 1781 -226 1815 -222
rect 1787 -232 1791 -226
rect 1706 -256 1739 -252
rect 1455 -275 1490 -271
rect 1120 -282 1124 -278
rect 1156 -281 1160 -278
rect 1107 -283 1124 -282
rect 1005 -288 1025 -284
rect 1041 -288 1056 -284
rect 1097 -286 1124 -283
rect 1005 -292 1009 -288
rect 1041 -291 1045 -288
rect 1097 -289 1103 -286
rect 992 -293 1009 -292
rect 847 -299 881 -295
rect 982 -296 1009 -293
rect 1138 -292 1142 -286
rect 853 -304 857 -299
rect 871 -304 875 -299
rect 895 -301 929 -297
rect 982 -299 988 -296
rect 901 -307 905 -301
rect 1023 -302 1027 -296
rect 1089 -300 1093 -294
rect 1107 -300 1111 -294
rect 1132 -295 1166 -292
rect 835 -325 854 -321
rect 862 -328 866 -314
rect 974 -310 978 -304
rect 992 -310 996 -304
rect 1017 -305 1051 -302
rect 1083 -303 1117 -300
rect 968 -313 1002 -310
rect 919 -325 923 -317
rect 1455 -315 1461 -275
rect 1498 -278 1502 -264
rect 1756 -258 1760 -245
rect 1805 -250 1809 -242
rect 1769 -254 1789 -250
rect 1805 -254 1817 -250
rect 1769 -258 1773 -254
rect 1805 -257 1809 -254
rect 1756 -259 1773 -258
rect 1746 -262 1773 -259
rect 1746 -265 1752 -262
rect 1787 -268 1791 -262
rect 1498 -279 1511 -278
rect 1520 -279 1539 -275
rect 1738 -276 1742 -270
rect 1756 -276 1760 -270
rect 1781 -271 1815 -268
rect 1498 -282 1523 -279
rect 1620 -280 1654 -276
rect 1732 -279 1766 -276
rect 1507 -283 1523 -282
rect 1537 -293 1541 -287
rect 1626 -288 1630 -280
rect 1489 -297 1493 -293
rect 1531 -296 1565 -293
rect 1483 -300 1517 -297
rect 1669 -289 1703 -285
rect 1675 -295 1679 -289
rect 1455 -321 1592 -315
rect 862 -329 875 -328
rect 884 -329 903 -325
rect 919 -329 956 -325
rect 862 -332 887 -329
rect 919 -332 923 -329
rect 871 -333 887 -332
rect 901 -343 905 -337
rect 853 -347 857 -343
rect 895 -346 929 -343
rect 1487 -346 1521 -342
rect 847 -350 881 -347
rect 1493 -351 1497 -346
rect 1511 -351 1515 -346
rect 1535 -348 1569 -344
rect 1584 -347 1592 -321
rect 1604 -319 1627 -315
rect 1604 -347 1610 -319
rect 1644 -321 1648 -308
rect 1657 -317 1677 -313
rect 1657 -321 1661 -317
rect 1644 -322 1661 -321
rect 1634 -325 1661 -322
rect 1634 -328 1640 -325
rect 1675 -331 1679 -325
rect 2244 -328 2248 -209
rect 2302 -212 2306 -198
rect 2302 -213 2315 -212
rect 2324 -213 2343 -209
rect 2302 -216 2327 -213
rect 2311 -217 2327 -216
rect 2341 -227 2345 -221
rect 2293 -231 2297 -227
rect 2335 -230 2369 -227
rect 2287 -234 2321 -231
rect 2560 -261 2564 -143
rect 2788 -217 2822 -213
rect 2603 -226 2637 -222
rect 2794 -225 2798 -217
rect 2609 -234 2613 -226
rect 2652 -235 2686 -231
rect 2658 -241 2662 -235
rect 2837 -226 2871 -222
rect 2843 -232 2847 -226
rect 2560 -265 2610 -261
rect 2627 -267 2631 -254
rect 2676 -259 2680 -251
rect 2722 -256 2795 -252
rect 2722 -259 2726 -256
rect 2812 -258 2816 -245
rect 2825 -254 2845 -250
rect 2825 -258 2829 -254
rect 2812 -259 2829 -258
rect 2640 -263 2660 -259
rect 2676 -263 2726 -259
rect 2802 -262 2829 -259
rect 2640 -267 2644 -263
rect 2676 -266 2680 -263
rect 2802 -265 2808 -262
rect 2627 -268 2644 -267
rect 2617 -271 2644 -268
rect 2843 -268 2847 -262
rect 2617 -274 2623 -271
rect 2658 -277 2662 -271
rect 2794 -276 2798 -270
rect 2812 -276 2816 -270
rect 2837 -271 2871 -268
rect 2609 -285 2613 -279
rect 2627 -285 2631 -279
rect 2652 -280 2686 -277
rect 2788 -279 2822 -276
rect 2603 -288 2637 -285
rect 2292 -306 2326 -302
rect 2298 -311 2302 -306
rect 2316 -311 2320 -306
rect 2340 -308 2374 -304
rect 2346 -314 2350 -308
rect 1626 -339 1630 -333
rect 1644 -339 1648 -333
rect 1669 -334 1703 -331
rect 2244 -332 2299 -328
rect 1620 -342 1654 -339
rect 1541 -354 1545 -348
rect 1464 -372 1494 -368
rect 1464 -398 1470 -372
rect 1502 -375 1506 -361
rect 1502 -376 1515 -375
rect 1524 -376 1543 -372
rect 1502 -379 1527 -376
rect 1511 -380 1527 -379
rect 1541 -390 1545 -384
rect 1493 -394 1497 -390
rect 1535 -393 1569 -390
rect 1487 -397 1521 -394
rect 2244 -456 2248 -332
rect 2307 -335 2311 -321
rect 2364 -332 2368 -324
rect 2307 -336 2320 -335
rect 2329 -336 2348 -332
rect 2364 -336 2387 -332
rect 2307 -339 2332 -336
rect 2364 -339 2368 -336
rect 2316 -340 2332 -339
rect 2346 -350 2350 -344
rect 2298 -354 2302 -350
rect 2340 -353 2374 -350
rect 2292 -357 2326 -354
rect 2384 -385 2387 -336
rect 2426 -350 2460 -346
rect 2432 -358 2436 -350
rect 2475 -359 2509 -355
rect 2481 -365 2485 -359
rect 2384 -389 2433 -385
rect 2450 -391 2454 -378
rect 2463 -387 2483 -383
rect 2463 -391 2467 -387
rect 2450 -392 2467 -391
rect 2440 -395 2467 -392
rect 2440 -398 2446 -395
rect 2481 -401 2485 -395
rect 2432 -409 2436 -403
rect 2450 -409 2454 -403
rect 2475 -404 2509 -401
rect 2426 -412 2460 -409
rect 2291 -434 2325 -430
rect 2297 -439 2301 -434
rect 2315 -439 2319 -434
rect 2339 -436 2373 -432
rect 2345 -442 2349 -436
rect 2244 -460 2298 -456
rect 2244 -489 2248 -460
rect 2306 -463 2310 -449
rect 2306 -464 2319 -463
rect 2328 -464 2347 -460
rect 2306 -467 2331 -464
rect 2315 -468 2331 -467
rect 2345 -478 2349 -472
rect 2297 -482 2301 -478
rect 2339 -481 2373 -478
rect 2291 -485 2325 -482
<< m2contact >>
rect 2266 -56 2271 -51
rect 2256 -87 2261 -82
rect 829 -217 834 -212
rect 950 -325 956 -320
<< metal2 >>
rect 2256 -82 2261 -42
rect 2271 -56 2329 -51
rect 2325 -82 2329 -56
rect 2315 -86 2329 -82
rect 880 -186 936 -182
rect 880 -212 884 -186
rect 817 -217 829 -212
rect 869 -216 884 -212
rect 468 -270 471 -263
rect 938 -287 943 -211
rect 1597 -217 1600 -138
rect 2441 -145 2444 -141
rect 2380 -148 2444 -145
rect 2228 -179 2328 -175
rect 2324 -205 2328 -179
rect 2314 -209 2328 -205
rect 2359 -210 2363 -201
rect 2380 -210 2383 -148
rect 2359 -213 2383 -210
rect 1630 -217 1633 -213
rect 2359 -216 2363 -213
rect 1574 -220 1633 -217
rect 1555 -276 1559 -267
rect 1574 -276 1578 -220
rect 1746 -256 1749 -252
rect 2861 -250 2865 -242
rect 2802 -256 2805 -252
rect 1097 -280 1100 -276
rect 1072 -283 1100 -280
rect 1555 -280 1578 -276
rect 1708 -259 1749 -256
rect 2749 -259 2805 -256
rect 2861 -254 2873 -250
rect 2861 -257 2865 -254
rect 1555 -282 1559 -280
rect 884 -291 943 -287
rect 982 -290 985 -286
rect 884 -321 888 -291
rect 874 -325 888 -321
rect 938 -352 943 -291
rect 950 -293 985 -290
rect 950 -313 956 -293
rect 1072 -308 1080 -283
rect 1693 -313 1697 -305
rect 1708 -313 1712 -259
rect 2617 -265 2620 -261
rect 2749 -263 2753 -259
rect 2588 -268 2620 -265
rect 2228 -302 2333 -297
rect 950 -320 956 -318
rect 1634 -319 1637 -315
rect 1610 -322 1637 -319
rect 1693 -317 1712 -313
rect 1693 -320 1697 -317
rect 1455 -341 1529 -337
rect 1525 -368 1529 -341
rect 1610 -347 1615 -322
rect 2329 -328 2333 -302
rect 2319 -332 2333 -328
rect 1514 -372 1529 -368
rect 1559 -372 1563 -364
rect 1559 -376 1580 -372
rect 1559 -379 1563 -376
rect 2499 -383 2503 -375
rect 2588 -383 2593 -268
rect 2440 -389 2443 -385
rect 2384 -392 2443 -389
rect 2499 -387 2593 -383
rect 2499 -390 2503 -387
rect 2228 -430 2332 -426
rect 2328 -456 2332 -430
rect 2318 -460 2332 -456
rect 2363 -461 2367 -452
rect 2384 -461 2387 -392
rect 2363 -464 2387 -461
rect 2363 -467 2367 -464
<< m3contact >>
rect 950 -318 956 -313
<< m123contact >>
rect 1817 -254 1822 -249
<< metal3 >>
rect 1455 -137 1526 -132
rect 1522 -165 1526 -137
rect 1511 -169 1526 -165
rect 914 -216 918 -208
rect 943 -216 947 -211
rect 914 -220 947 -216
rect 914 -223 918 -220
rect 377 -263 386 -259
rect 943 -286 947 -220
rect 1455 -244 1523 -239
rect 1518 -271 1523 -244
rect 1817 -249 1822 -138
rect 1510 -275 1523 -271
rect 943 -290 975 -286
rect 956 -318 1038 -313
<< labels >>
rlabel polycontact 975 -290 979 -286 1 p1g0
rlabel polycontact 898 -220 902 -216 1 p1g0n
rlabel pdcontact 914 -208 918 -198 1 p1g0
rlabel ndcontact 914 -228 918 -223 1 p1g0
rlabel polycontact 870 -325 874 -321 1 p1
rlabel polycontact 865 -216 869 -212 1 p1
rlabel polycontact 1090 -280 1094 -276 1 or1c2
rlabel metal1 1052 -288 1056 -276 1 or1c2
rlabel ndcontact 1041 -296 1045 -291 1 or1c2
rlabel pdcontact 1041 -276 1045 -266 1 or1c2
rlabel polycontact 1025 -288 1029 -284 1 or1c2n
rlabel metal1 997 -296 1009 -292 1 or1c2n
rlabel ndcontact 982 -304 988 -299 1 or1c2n
rlabel pdcontact 992 -279 996 -259 1 or1c2n
rlabel polycontact 854 -325 858 -321 1 p0c0
rlabel ndiffusion 856 -234 862 -224 1 and2nmc2
rlabel ndiffusion 861 -343 867 -333 1 and1nmc2
rlabel metal1 879 -333 887 -329 1 p1p0c0n
rlabel pdcontact 862 -314 866 -304 1 p1p0c0n
rlabel ndcontact 871 -343 875 -333 1 p1p0c0n
rlabel polycontact 903 -329 907 -325 1 p1p0c0n
rlabel metal1 923 -329 932 -325 1 p1p0c0
rlabel pdcontact 919 -317 923 -307 1 p1p0c0
rlabel ndcontact 919 -337 923 -332 1 p1p0c0
rlabel polycontact 985 -290 989 -286 1 p1p0c0
rlabel metal3 914 -220 926 -216 1 p1g0
rlabel ndcontact 866 -234 870 -224 1 p1g0n
rlabel pdcontact 857 -205 861 -195 1 p1g0n
rlabel polycontact 849 -217 853 -212 1 g0
rlabel pdiffusion 982 -279 988 -259 1 or1pmc2
rlabel pdiffusion 1097 -269 1103 -249 1 or2pmc2
rlabel pdcontact 1107 -269 1111 -249 1 c2n
rlabel ndcontact 1097 -294 1103 -289 1 c2n
rlabel polycontact 1140 -278 1144 -274 1 c2n
rlabel metal1 1170 -278 1182 -274 1 c2
rlabel pdcontact 1156 -266 1160 -256 1 c2
rlabel ndcontact 1156 -286 1160 -281 1 c2
rlabel polycontact 1100 -280 1104 -276 1 g1
rlabel pdcontact 1089 -269 1093 -249 1 vdd
rlabel pdcontact 974 -279 978 -259 1 vdd
rlabel pdcontact 896 -208 900 -198 1 vdd
rlabel pdcontact 866 -205 870 -195 1 vdd
rlabel pdcontact 848 -205 852 -195 1 vdd
rlabel pdcontact 871 -314 875 -304 1 vdd
rlabel pdcontact 853 -314 857 -304 1 vdd
rlabel pdcontact 901 -317 905 -307 1 vdd
rlabel pdcontact 1023 -276 1027 -266 1 vdd
rlabel pdcontact 1138 -266 1142 -256 1 vdd
rlabel ndcontact 1138 -286 1142 -281 1 gnd
rlabel ndcontact 1107 -294 1111 -289 1 gnd
rlabel ndcontact 1089 -294 1093 -289 1 gnd
rlabel ndcontact 1023 -296 1027 -291 1 gnd
rlabel ndcontact 992 -304 996 -299 1 gnd
rlabel ndcontact 974 -304 978 -299 1 gnd
rlabel ndcontact 901 -337 905 -332 1 gnd
rlabel ndcontact 896 -228 900 -223 1 gnd
rlabel ndcontact 848 -234 852 -224 1 gnd
rlabel ndcontact 853 -343 857 -333 1 gnd
rlabel metal1 890 -237 924 -234 1 gnd
rlabel metal1 842 -241 876 -238 1 gnd
rlabel metal1 847 -350 881 -347 1 gnd
rlabel metal1 895 -346 929 -343 1 gnd
rlabel metal1 968 -313 1002 -310 1 gnd
rlabel metal1 1017 -305 1051 -302 1 gnd
rlabel metal1 1083 -303 1117 -300 1 gnd
rlabel metal1 1132 -295 1166 -292 1 gnd
rlabel metal1 1132 -250 1166 -246 1 vdd
rlabel metal1 1083 -241 1117 -237 1 vdd
rlabel metal1 1017 -260 1051 -256 1 vdd
rlabel metal1 968 -251 1002 -247 1 vdd
rlabel metal1 895 -301 929 -297 1 vdd
rlabel metal1 847 -299 881 -295 1 vdd
rlabel metal1 890 -192 924 -188 1 vdd
rlabel metal1 842 -190 876 -186 1 vdd
rlabel polysilicon 1104 -280 1106 -276 1 g1
rlabel pdcontact 1693 -305 1697 -295 1 or2c3
rlabel ndcontact 1693 -325 1697 -320 1 or2c3
rlabel polycontact 1507 -169 1511 -165 1 p1g0
rlabel pdcontact 1555 -267 1559 -257 1 p2p1p0c0
rlabel ndcontact 1555 -287 1559 -282 1 p2p1p0c0
rlabel polycontact 1506 -275 1510 -271 1 p1p0c0
rlabel polycontact 1673 -215 1677 -211 1 orc3n
rlabel metal1 1647 -223 1657 -219 1 orc3n
rlabel ndcontact 1630 -231 1636 -226 1 orc3n
rlabel pdcontact 1640 -206 1644 -186 1 orc3n
rlabel pdcontact 1644 -308 1648 -288 1 or2c3n
rlabel ndcontact 1634 -333 1640 -328 1 or2c3n
rlabel metal1 1648 -325 1657 -321 1 or2c3n
rlabel polycontact 1677 -317 1681 -313 1 or2c3n
rlabel metal2 1699 -317 1708 -313 1 or2c3
rlabel polycontact 1749 -256 1753 -252 1 or2c3
rlabel polycontact 1739 -256 1743 -252 1 orc3
rlabel metal1 1696 -215 1706 -211 1 orc3
rlabel ndcontact 1689 -223 1693 -218 1 orc3
rlabel pdcontact 1689 -203 1693 -193 1 orc3
rlabel metal1 1812 -254 1817 -250 1 c3
rlabel metal3 1817 -254 1822 -243 1 c3
rlabel ndcontact 1805 -262 1809 -257 1 c3
rlabel pdcontact 1805 -242 1809 -232 1 c3
rlabel polycontact 1789 -254 1793 -250 1 c3n
rlabel metal1 1769 -262 1773 -250 1 c3n
rlabel ndcontact 1746 -270 1752 -265 1 c3n
rlabel pdcontact 1756 -245 1760 -225 1 c3n
rlabel pdiffusion 1746 -245 1752 -225 1 or1pmc3
rlabel pdiffusion 1634 -308 1640 -288 1 or2pmc3
rlabel polycontact 1637 -319 1641 -315 1 p2g1
rlabel polycontact 1627 -319 1631 -315 1 g2
rlabel pdiffusion 1630 -206 1636 -186 1 or3pmc3
rlabel polycontact 1623 -217 1627 -213 1 p2p1g0
rlabel polycontact 1633 -217 1637 -213 1 p2p1p0c0
rlabel ndiffusion 1498 -187 1504 -177 1 and3nmc3
rlabel metal1 1560 -173 1572 -169 1 p2p1g0
rlabel ndcontact 1556 -181 1560 -176 1 p2p1g0
rlabel pdcontact 1556 -161 1560 -151 1 p2p1g0
rlabel polycontact 1540 -173 1544 -169 1 p2p1g0n
rlabel ndcontact 1508 -187 1512 -177 1 p2p1g0n
rlabel pdcontact 1499 -158 1503 -148 1 p2p1g0n
rlabel metal2 1563 -376 1574 -372 1 p2g1
rlabel polycontact 1543 -376 1547 -372 1 p2g1n
rlabel metal1 1519 -380 1527 -376 1 p2g1n
rlabel ndcontact 1511 -390 1515 -380 1 p2g1n
rlabel pdcontact 1502 -361 1506 -351 1 p2g1n
rlabel ndiffusion 1501 -390 1507 -380 1 and1nmc3
rlabel ndiffusion 1497 -293 1503 -283 1 and2nmc3
rlabel metal2 1561 -280 1571 -276 1 p2p1p0c0
rlabel polycontact 1539 -279 1543 -275 1 p2p1p0c0n
rlabel ndcontact 1507 -293 1511 -283 1 p2p1p0c0n
rlabel pdcontact 1498 -264 1502 -254 1 p2p1p0c0n
rlabel polycontact 1491 -169 1495 -165 1 p2
rlabel polycontact 1490 -275 1494 -271 1 p2
rlabel polycontact 1494 -372 1498 -368 1 p2
rlabel pdcontact 1538 -161 1542 -151 1 vdd
rlabel pdcontact 1508 -158 1512 -148 1 vdd
rlabel pdcontact 1490 -158 1494 -148 1 vdd
rlabel pdcontact 1507 -264 1511 -254 1 vdd
rlabel pdcontact 1489 -264 1493 -254 1 vdd
rlabel pdcontact 1511 -361 1515 -351 1 vdd
rlabel pdcontact 1493 -361 1497 -351 1 vdd
rlabel pdcontact 1541 -364 1545 -354 1 vdd
rlabel pdcontact 1537 -267 1541 -257 1 vdd
rlabel pdcontact 1675 -305 1679 -295 1 vdd
rlabel pdcontact 1671 -203 1675 -193 1 vdd
rlabel pdcontact 1622 -206 1626 -186 1 vdd
rlabel pdcontact 1626 -308 1630 -288 1 vdd
rlabel pdcontact 1738 -245 1742 -225 1 vdd
rlabel pdcontact 1787 -242 1791 -232 1 vdd
rlabel ndcontact 1787 -262 1791 -257 1 gnd
rlabel ndcontact 1756 -270 1760 -265 1 gnd
rlabel ndcontact 1738 -270 1742 -265 1 gnd
rlabel ndcontact 1675 -325 1679 -320 1 gnd
rlabel ndcontact 1671 -223 1675 -218 1 gnd
rlabel ndcontact 1640 -231 1644 -226 1 gnd
rlabel ndcontact 1622 -231 1626 -226 1 gnd
rlabel ndcontact 1644 -333 1648 -328 1 gnd
rlabel ndcontact 1626 -333 1630 -328 1 gnd
rlabel ndcontact 1541 -384 1545 -379 1 gnd
rlabel ndcontact 1537 -287 1541 -282 1 gnd
rlabel ndcontact 1538 -181 1542 -176 1 gnd
rlabel ndcontact 1490 -187 1494 -177 1 gnd
rlabel ndcontact 1489 -293 1493 -283 1 gnd
rlabel ndcontact 1493 -390 1497 -380 1 gnd
rlabel metal1 1535 -393 1569 -390 1 gnd
rlabel metal1 1487 -397 1521 -394 1 gnd
rlabel metal1 1532 -190 1566 -187 1 gnd
rlabel metal1 1484 -194 1518 -191 1 gnd
rlabel metal1 1483 -300 1517 -297 1 gnd
rlabel metal1 1531 -296 1565 -293 1 gnd
rlabel metal1 1669 -334 1703 -331 1 gnd
rlabel metal1 1620 -342 1654 -339 1 gnd
rlabel metal1 1665 -232 1699 -229 1 gnd
rlabel metal1 1616 -240 1650 -237 1 gnd
rlabel metal1 1732 -279 1766 -276 1 gnd
rlabel metal1 1781 -271 1815 -268 1 gnd
rlabel metal1 1781 -226 1815 -222 1 vdd
rlabel metal1 1732 -217 1766 -213 1 vdd
rlabel metal1 1669 -289 1703 -285 1 vdd
rlabel metal1 1620 -280 1654 -276 1 vdd
rlabel metal1 1665 -187 1699 -183 1 vdd
rlabel metal1 1616 -178 1650 -174 1 vdd
rlabel metal1 1535 -348 1569 -344 1 vdd
rlabel metal1 1487 -346 1521 -342 1 vdd
rlabel metal1 1531 -251 1565 -247 1 vdd
rlabel metal1 1483 -249 1517 -245 1 vdd
rlabel metal1 1532 -145 1566 -141 1 vdd
rlabel metal1 1484 -143 1518 -139 1 vdd
rlabel pdcontact 1559 -364 1563 -354 1 p2g1
rlabel ndcontact 1559 -384 1563 -379 1 p2g1
rlabel polycontact 1510 -372 1514 -368 1 g1
rlabel polysilicon 1508 -372 1510 -368 1 g1
rlabel metal2 2868 -254 2873 -250 1 c4
rlabel pdcontact 2861 -242 2865 -232 1 c4
rlabel ndcontact 2861 -262 2865 -257 1 c4
rlabel pdcontact 2499 -375 2503 -365 1 or2c4
rlabel ndcontact 2499 -395 2503 -390 1 or2c4
rlabel polycontact 2311 -86 2315 -82 1 p2p1g0
rlabel pdcontact 2359 -201 2363 -191 1 p3p2p1p0c0
rlabel ndcontact 2359 -221 2363 -216 1 p3p2p1p0c0
rlabel polycontact 2310 -209 2314 -205 1 p2p1p0c0
rlabel pdcontact 2363 -452 2367 -442 1 p3p2g1
rlabel ndcontact 2363 -472 2367 -467 1 p3p2g1
rlabel polycontact 2314 -460 2318 -456 1 p2g1
rlabel pdcontact 2346 -324 2350 -314 1 vdd
rlabel ndcontact 2843 -262 2847 -257 1 gnd
rlabel ndcontact 2812 -270 2816 -265 1 gnd
rlabel ndcontact 2794 -270 2798 -265 1 gnd
rlabel pdcontact 2843 -242 2847 -232 1 vdd
rlabel pdcontact 2794 -245 2798 -225 1 vdd
rlabel polycontact 2845 -254 2849 -250 1 coutn
rlabel metal1 2817 -262 2822 -258 1 coutn
rlabel ndcontact 2802 -270 2808 -265 1 coutn
rlabel pdcontact 2812 -245 2816 -225 1 coutn
rlabel pdiffusion 2802 -245 2808 -225 1 or0pmc4
rlabel polycontact 2795 -256 2799 -252 1 or1c4
rlabel metal1 2686 -263 2694 -259 1 or1c4
rlabel ndcontact 2676 -271 2680 -266 1 or1c4
rlabel pdcontact 2676 -251 2680 -241 1 or1c4
rlabel polycontact 2660 -263 2664 -259 1 or1c4n
rlabel metal1 2638 -271 2642 -267 1 or1c4n
rlabel ndcontact 2617 -279 2623 -274 1 or1c4n
rlabel pdcontact 2627 -254 2631 -234 1 or1c4n
rlabel ndcontact 2658 -271 2662 -266 1 gnd
rlabel ndcontact 2627 -279 2631 -274 1 gnd
rlabel ndcontact 2609 -279 2613 -274 1 gnd
rlabel pdcontact 2658 -251 2662 -241 1 vdd
rlabel pdcontact 2609 -254 2613 -234 1 vdd
rlabel pdiffusion 2617 -254 2623 -234 1 or1pmc4
rlabel polycontact 2620 -265 2624 -261 1 or2c4
rlabel metal2 2523 -387 2531 -383 1 or2c4
rlabel polycontact 2483 -387 2487 -383 1 or2c4n
rlabel metal1 2457 -395 2463 -391 1 or2c4n
rlabel ndcontact 2440 -403 2446 -398 1 or2c4n
rlabel pdcontact 2450 -378 2454 -358 1 or2c4n
rlabel pdiffusion 2440 -378 2446 -358 1 or2pmc4
rlabel ndcontact 2481 -395 2485 -390 1 gnd
rlabel ndcontact 2450 -403 2454 -398 1 gnd
rlabel ndcontact 2432 -403 2436 -398 1 gnd
rlabel pdcontact 2481 -375 2485 -365 1 vdd
rlabel pdcontact 2432 -378 2436 -358 1 vdd
rlabel polycontact 2610 -265 2614 -261 1 or3c4
rlabel metal1 2509 -143 2514 -139 1 or3c4
rlabel ndcontact 2500 -151 2504 -146 1 or3c4
rlabel pdcontact 2500 -131 2504 -121 1 or3c4
rlabel polycontact 2484 -143 2488 -139 1 or3nc4
rlabel metal1 2464 -151 2468 -143 1 or3nc4
rlabel ndcontact 2441 -159 2447 -154 1 or3nc4
rlabel pdcontact 2451 -134 2455 -114 1 or3nc4
rlabel pdiffusion 2441 -134 2447 -114 1 or3pmc4
rlabel ndcontact 2482 -151 2486 -146 1 gnd
rlabel ndcontact 2451 -159 2455 -154 1 gnd
rlabel ndcontact 2433 -159 2437 -154 1 gnd
rlabel pdcontact 2482 -131 2486 -121 1 vdd
rlabel pdcontact 2433 -134 2437 -114 1 vdd
rlabel polycontact 2434 -145 2438 -141 1 p3p2p1g0
rlabel ndcontact 2346 -344 2350 -339 1 gnd
rlabel pdcontact 2345 -452 2349 -442 1 vdd
rlabel ndcontact 2345 -472 2349 -467 1 gnd
rlabel ndcontact 2297 -478 2301 -468 1 gnd
rlabel pdcontact 2315 -449 2319 -439 1 vdd
rlabel pdcontact 2297 -449 2301 -439 1 vdd
rlabel polycontact 2295 -87 2299 -82 1 p3
rlabel metal1 2373 -90 2383 -86 1 p3p2p1g0
rlabel pdcontact 2360 -78 2364 -68 1 p3p2p1g0
rlabel ndcontact 2360 -98 2364 -93 1 p3p2p1g0
rlabel ndcontact 2342 -98 2346 -93 1 gnd
rlabel ndiffusion 2302 -104 2308 -94 1 and4nmc4
rlabel polycontact 2344 -90 2348 -86 1 p3p2p1g0n
rlabel metal1 2318 -94 2328 -90 1 p3p2p1g0n
rlabel ndcontact 2312 -104 2316 -94 1 p3p2p1g0n
rlabel pdcontact 2303 -75 2307 -65 1 p3p2p1g0n
rlabel pdcontact 2342 -78 2346 -68 1 vdd
rlabel pdcontact 2312 -75 2316 -65 1 vdd
rlabel pdcontact 2294 -75 2298 -65 1 vdd
rlabel ndcontact 2294 -104 2298 -94 1 gnd
rlabel ndcontact 2293 -227 2297 -217 1 gnd
rlabel ndcontact 2341 -221 2345 -216 1 gnd
rlabel polycontact 2444 -145 2448 -141 1 p3p2p1p0c0
rlabel metal2 2369 -213 2380 -210 1 p3p2p1p0c0
rlabel polycontact 2343 -213 2347 -209 1 p3p2p1p0c0n
rlabel ndiffusion 2301 -227 2307 -217 1 and3nmc4
rlabel ndcontact 2311 -227 2315 -217 1 p3p2p1p0c0n
rlabel pdcontact 2302 -198 2306 -188 1 p3p2p1p0c0n
rlabel pdcontact 2311 -198 2315 -188 1 vdd
rlabel pdcontact 2293 -198 2297 -188 1 vdd
rlabel pdcontact 2341 -201 2345 -191 1 vdd
rlabel polycontact 2433 -389 2437 -385 1 p3g2
rlabel metal1 2377 -336 2384 -332 1 p3g2
rlabel ndcontact 2364 -344 2368 -339 1 p3g2
rlabel pdcontact 2364 -324 2368 -314 1 p3g2
rlabel polycontact 2348 -336 2352 -332 1 p3g2n
rlabel metal1 2324 -340 2332 -336 1 p3g2n
rlabel ndcontact 2316 -350 2320 -340 1 p3g2n
rlabel pdcontact 2307 -321 2311 -311 1 p3g2n
rlabel pdcontact 2316 -321 2320 -311 1 vdd
rlabel pdcontact 2298 -321 2302 -311 1 vdd
rlabel ndcontact 2298 -350 2302 -340 1 gnd
rlabel ndiffusion 2306 -350 2312 -340 1 and2nmc4
rlabel ndiffusion 2305 -478 2311 -468 1 and1nmc4
rlabel metal2 2375 -464 2384 -461 1 p2p3g1
rlabel polycontact 2347 -464 2351 -460 1 p2p3g1n
rlabel ndcontact 2315 -478 2319 -468 1 p2p3g1n
rlabel pdcontact 2306 -449 2310 -439 1 p2p3g1n
rlabel polycontact 2805 -256 2809 -252 1 g3
rlabel polycontact 2294 -209 2298 -205 1 p3
rlabel polycontact 2299 -332 2303 -328 1 p3
rlabel polycontact 2298 -460 2302 -456 1 p3
rlabel metal1 2339 -481 2373 -478 1 gnd
rlabel metal1 2291 -485 2325 -482 1 gnd
rlabel metal1 2340 -353 2374 -350 1 gnd
rlabel metal1 2292 -357 2326 -354 1 gnd
rlabel metal1 2335 -230 2369 -227 1 gnd
rlabel metal1 2287 -234 2321 -231 1 gnd
rlabel metal1 2336 -107 2370 -104 1 gnd
rlabel metal1 2288 -111 2322 -108 1 gnd
rlabel metal1 2476 -160 2510 -157 1 gnd
rlabel metal1 2427 -168 2461 -165 1 gnd
rlabel metal1 2475 -404 2509 -401 1 gnd
rlabel metal1 2426 -412 2460 -409 1 gnd
rlabel metal1 2603 -288 2637 -285 1 gnd
rlabel metal1 2652 -280 2686 -277 1 gnd
rlabel metal1 2788 -279 2822 -276 1 gnd
rlabel metal1 2837 -271 2871 -268 1 gnd
rlabel metal1 2837 -226 2871 -222 1 vdd
rlabel metal1 2788 -217 2822 -213 1 vdd
rlabel metal1 2652 -235 2686 -231 1 vdd
rlabel metal1 2603 -226 2637 -222 1 vdd
rlabel metal1 2476 -115 2510 -111 1 vdd
rlabel metal1 2427 -106 2461 -102 1 vdd
rlabel metal1 2336 -62 2370 -58 1 vdd
rlabel metal1 2288 -60 2322 -56 1 vdd
rlabel metal1 2335 -185 2369 -181 1 vdd
rlabel metal1 2287 -183 2321 -179 1 vdd
rlabel metal1 2475 -359 2509 -355 1 vdd
rlabel metal1 2426 -350 2460 -346 1 vdd
rlabel metal1 2339 -436 2373 -432 1 vdd
rlabel metal1 2291 -434 2325 -430 1 vdd
rlabel metal1 2340 -308 2374 -304 1 vdd
rlabel metal1 2292 -306 2326 -302 1 vdd
rlabel polycontact 2315 -332 2319 -328 1 g2
rlabel polysilicon 2313 -332 2315 -328 1 g2
rlabel polysilicon 2809 -256 2811 -252 1 g3
rlabel polysilicon 2448 -145 2450 -141 1 p3p2p1p0c0
rlabel polycontact 2443 -389 2447 -385 1 p3p2g1
rlabel polysilicon 2447 -389 2449 -385 1 p3p2g1
rlabel polycontact 461 -267 465 -263 1 p0c0
rlabel metal1 426 -267 435 -263 1 p0c0
rlabel ndcontact 422 -275 426 -270 1 p0c0
rlabel pdcontact 422 -255 426 -245 1 p0c0
rlabel polycontact 406 -267 410 -263 1 p0c0n
rlabel metal1 380 -271 390 -267 1 p0c0n
rlabel ndcontact 374 -281 378 -271 1 p0c0n
rlabel pdcontact 365 -252 369 -242 1 p0c0n
rlabel ndiffusion 364 -281 370 -271 1 andnmc1
rlabel ndcontact 527 -273 531 -268 1 c1
rlabel pdcontact 527 -253 531 -243 1 c1
rlabel polycontact 511 -265 515 -261 1 c1n
rlabel ndcontact 468 -281 474 -276 1 c1n
rlabel pdcontact 478 -256 482 -236 1 c1n
rlabel pdiffusion 468 -256 474 -236 1 orpmc1
rlabel polycontact 471 -267 475 -263 1 g0
rlabel polycontact 357 -263 361 -259 1 p0
rlabel pdcontact 460 -256 464 -236 1 vdd
rlabel pdcontact 509 -253 513 -243 1 vdd
rlabel pdcontact 404 -255 408 -245 1 vdd
rlabel pdcontact 374 -252 378 -242 1 vdd
rlabel pdcontact 356 -252 360 -242 1 vdd
rlabel ndcontact 509 -273 513 -268 1 gnd
rlabel ndcontact 478 -281 482 -276 1 gnd
rlabel ndcontact 460 -281 464 -276 1 gnd
rlabel ndcontact 404 -275 408 -270 1 gnd
rlabel ndcontact 356 -281 360 -271 1 gnd
rlabel metal1 350 -288 384 -285 1 gnd
rlabel metal1 398 -284 432 -281 1 gnd
rlabel metal1 454 -290 488 -287 1 gnd
rlabel metal1 503 -282 537 -279 1 gnd
rlabel metal1 503 -237 537 -233 1 vdd
rlabel metal1 454 -228 488 -224 1 vdd
rlabel metal1 398 -239 432 -235 1 vdd
rlabel metal1 350 -237 384 -233 1 vdd
rlabel polycontact 373 -263 377 -259 1 c0
rlabel polysilicon 475 -267 477 -263 1 g0
rlabel polysilicon 371 -263 373 -259 1 c0
<< end >>
