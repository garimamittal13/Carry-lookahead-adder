magic
tech scmos
timestamp 1732093082
<< error_p >>
rect 877 -1178 879 -1173
<< nwell >>
rect -353 -1133 -319 -1107
rect -307 -1123 -273 -1098
rect -259 -1126 -225 -1100
rect -353 -1189 -319 -1163
rect -305 -1189 -271 -1164
rect -257 -1192 -223 -1166
rect -199 -1169 -165 -1131
rect -150 -1166 -116 -1140
rect 82 -1150 116 -1124
rect 128 -1140 162 -1115
rect 176 -1143 210 -1117
rect 587 -1139 621 -1113
rect 633 -1129 667 -1104
rect 681 -1132 715 -1106
rect 1043 -1126 1077 -1100
rect 1089 -1116 1123 -1091
rect 1137 -1119 1171 -1093
rect 82 -1206 116 -1180
rect 130 -1206 164 -1181
rect 178 -1209 212 -1183
rect 236 -1186 270 -1148
rect 285 -1183 319 -1157
rect 587 -1195 621 -1169
rect 635 -1195 669 -1170
rect 683 -1198 717 -1172
rect 741 -1175 775 -1137
rect 790 -1172 824 -1146
rect 1043 -1182 1077 -1156
rect 1091 -1182 1125 -1157
rect 1139 -1185 1173 -1159
rect 1197 -1162 1231 -1124
rect 1246 -1159 1280 -1133
rect -337 -1298 -303 -1273
rect -289 -1301 -255 -1275
rect 133 -1297 167 -1272
rect 181 -1300 215 -1274
rect 627 -1285 661 -1260
rect 1078 -1261 1112 -1236
rect 675 -1288 709 -1262
rect 1126 -1264 1160 -1238
<< ntransistor >>
rect -341 -1147 -339 -1142
rect -296 -1146 -294 -1136
rect -286 -1146 -284 -1136
rect -247 -1140 -245 -1135
rect 1055 -1140 1057 -1135
rect 1100 -1139 1102 -1129
rect 1110 -1139 1112 -1129
rect 1149 -1133 1151 -1128
rect -341 -1203 -339 -1198
rect 94 -1164 96 -1159
rect 139 -1163 141 -1153
rect 149 -1163 151 -1153
rect 188 -1157 190 -1152
rect 599 -1153 601 -1148
rect 644 -1152 646 -1142
rect 654 -1152 656 -1142
rect 693 -1146 695 -1141
rect -138 -1180 -136 -1175
rect -188 -1188 -186 -1183
rect -178 -1188 -176 -1183
rect -294 -1212 -292 -1202
rect -284 -1212 -282 -1202
rect -245 -1206 -243 -1201
rect 94 -1220 96 -1215
rect 297 -1197 299 -1192
rect 247 -1205 249 -1200
rect 257 -1205 259 -1200
rect 599 -1209 601 -1204
rect 802 -1186 804 -1181
rect 752 -1194 754 -1189
rect 762 -1194 764 -1189
rect 1055 -1196 1057 -1191
rect 1258 -1173 1260 -1168
rect 1208 -1181 1210 -1176
rect 1218 -1181 1220 -1176
rect 1102 -1205 1104 -1195
rect 1112 -1205 1114 -1195
rect 1151 -1199 1153 -1194
rect 646 -1218 648 -1208
rect 656 -1218 658 -1208
rect 695 -1212 697 -1207
rect 141 -1229 143 -1219
rect 151 -1229 153 -1219
rect 190 -1223 192 -1218
rect 1089 -1284 1091 -1274
rect 1099 -1284 1101 -1274
rect 1138 -1278 1140 -1273
rect 638 -1308 640 -1298
rect 648 -1308 650 -1298
rect 687 -1302 689 -1297
rect -326 -1321 -324 -1311
rect -316 -1321 -314 -1311
rect -277 -1315 -275 -1310
rect 144 -1320 146 -1310
rect 154 -1320 156 -1310
rect 193 -1314 195 -1309
<< ptransistor >>
rect -296 -1117 -294 -1107
rect -286 -1117 -284 -1107
rect 1100 -1110 1102 -1100
rect 1110 -1110 1112 -1100
rect -341 -1127 -339 -1117
rect -247 -1120 -245 -1110
rect 644 -1123 646 -1113
rect 654 -1123 656 -1113
rect 139 -1134 141 -1124
rect 149 -1134 151 -1124
rect -188 -1163 -186 -1143
rect -178 -1163 -176 -1143
rect 94 -1144 96 -1134
rect -138 -1160 -136 -1150
rect 188 -1137 190 -1127
rect 599 -1133 601 -1123
rect 693 -1126 695 -1116
rect 1055 -1120 1057 -1110
rect 1149 -1113 1151 -1103
rect -341 -1183 -339 -1173
rect -294 -1183 -292 -1173
rect -284 -1183 -282 -1173
rect -245 -1186 -243 -1176
rect 247 -1180 249 -1160
rect 257 -1180 259 -1160
rect 297 -1177 299 -1167
rect 752 -1169 754 -1149
rect 762 -1169 764 -1149
rect 1208 -1156 1210 -1136
rect 1218 -1156 1220 -1136
rect 1258 -1153 1260 -1143
rect 802 -1166 804 -1156
rect 94 -1200 96 -1190
rect 141 -1200 143 -1190
rect 151 -1200 153 -1190
rect 190 -1203 192 -1193
rect 599 -1189 601 -1179
rect 646 -1189 648 -1179
rect 656 -1189 658 -1179
rect 695 -1192 697 -1182
rect 1055 -1176 1057 -1166
rect 1102 -1176 1104 -1166
rect 1112 -1176 1114 -1166
rect 1151 -1179 1153 -1169
rect 1089 -1255 1091 -1245
rect 1099 -1255 1101 -1245
rect 638 -1279 640 -1269
rect 648 -1279 650 -1269
rect -326 -1292 -324 -1282
rect -316 -1292 -314 -1282
rect -277 -1295 -275 -1285
rect 144 -1291 146 -1281
rect 154 -1291 156 -1281
rect 193 -1294 195 -1284
rect 687 -1282 689 -1272
rect 1138 -1258 1140 -1248
<< ndiffusion >>
rect -343 -1147 -341 -1142
rect -339 -1147 -329 -1142
rect -297 -1146 -296 -1136
rect -294 -1146 -286 -1136
rect -284 -1146 -283 -1136
rect -249 -1140 -247 -1135
rect -245 -1140 -235 -1135
rect 1053 -1140 1055 -1135
rect 1057 -1140 1067 -1135
rect 1099 -1139 1100 -1129
rect 1102 -1139 1110 -1129
rect 1112 -1139 1113 -1129
rect 1147 -1133 1149 -1128
rect 1151 -1133 1161 -1128
rect -343 -1203 -341 -1198
rect -339 -1203 -329 -1198
rect 92 -1164 94 -1159
rect 96 -1164 106 -1159
rect 138 -1163 139 -1153
rect 141 -1163 149 -1153
rect 151 -1163 152 -1153
rect 186 -1157 188 -1152
rect 190 -1157 200 -1152
rect 597 -1153 599 -1148
rect 601 -1153 611 -1148
rect 643 -1152 644 -1142
rect 646 -1152 654 -1142
rect 656 -1152 657 -1142
rect 691 -1146 693 -1141
rect 695 -1146 705 -1141
rect -140 -1180 -138 -1175
rect -136 -1180 -126 -1175
rect -189 -1188 -188 -1183
rect -186 -1188 -185 -1183
rect -179 -1188 -178 -1183
rect -176 -1188 -175 -1183
rect -295 -1212 -294 -1202
rect -292 -1212 -284 -1202
rect -282 -1212 -281 -1202
rect -247 -1206 -245 -1201
rect -243 -1206 -233 -1201
rect 92 -1220 94 -1215
rect 96 -1220 106 -1215
rect 295 -1197 297 -1192
rect 299 -1197 309 -1192
rect 246 -1205 247 -1200
rect 249 -1205 250 -1200
rect 256 -1205 257 -1200
rect 259 -1205 260 -1200
rect 597 -1209 599 -1204
rect 601 -1209 611 -1204
rect 800 -1186 802 -1181
rect 804 -1186 814 -1181
rect 751 -1194 752 -1189
rect 754 -1194 755 -1189
rect 761 -1194 762 -1189
rect 764 -1194 765 -1189
rect 1053 -1196 1055 -1191
rect 1057 -1196 1067 -1191
rect 1256 -1173 1258 -1168
rect 1260 -1173 1270 -1168
rect 1207 -1181 1208 -1176
rect 1210 -1181 1211 -1176
rect 1217 -1181 1218 -1176
rect 1220 -1181 1221 -1176
rect 1101 -1205 1102 -1195
rect 1104 -1205 1112 -1195
rect 1114 -1205 1115 -1195
rect 1149 -1199 1151 -1194
rect 1153 -1199 1163 -1194
rect 645 -1218 646 -1208
rect 648 -1218 656 -1208
rect 658 -1218 659 -1208
rect 693 -1212 695 -1207
rect 697 -1212 707 -1207
rect 140 -1229 141 -1219
rect 143 -1229 151 -1219
rect 153 -1229 154 -1219
rect 188 -1223 190 -1218
rect 192 -1223 202 -1218
rect 1088 -1284 1089 -1274
rect 1091 -1284 1099 -1274
rect 1101 -1284 1102 -1274
rect 1136 -1278 1138 -1273
rect 1140 -1278 1150 -1273
rect 637 -1308 638 -1298
rect 640 -1308 648 -1298
rect 650 -1308 651 -1298
rect 685 -1302 687 -1297
rect 689 -1302 699 -1297
rect -327 -1321 -326 -1311
rect -324 -1321 -316 -1311
rect -314 -1321 -313 -1311
rect -279 -1315 -277 -1310
rect -275 -1315 -265 -1310
rect 143 -1320 144 -1310
rect 146 -1320 154 -1310
rect 156 -1320 157 -1310
rect 191 -1314 193 -1309
rect 195 -1314 205 -1309
<< pdiffusion >>
rect -297 -1117 -296 -1107
rect -294 -1117 -292 -1107
rect -288 -1117 -286 -1107
rect -284 -1117 -283 -1107
rect 1099 -1110 1100 -1100
rect 1102 -1110 1104 -1100
rect 1108 -1110 1110 -1100
rect 1112 -1110 1113 -1100
rect -343 -1127 -341 -1117
rect -339 -1127 -329 -1117
rect -249 -1120 -247 -1110
rect -245 -1120 -235 -1110
rect 643 -1123 644 -1113
rect 646 -1123 648 -1113
rect 652 -1123 654 -1113
rect 656 -1123 657 -1113
rect 138 -1134 139 -1124
rect 141 -1134 143 -1124
rect 147 -1134 149 -1124
rect 151 -1134 152 -1124
rect -189 -1163 -188 -1143
rect -186 -1163 -178 -1143
rect -176 -1163 -175 -1143
rect 92 -1144 94 -1134
rect 96 -1144 106 -1134
rect -140 -1160 -138 -1150
rect -136 -1160 -126 -1150
rect 186 -1137 188 -1127
rect 190 -1137 200 -1127
rect 597 -1133 599 -1123
rect 601 -1133 611 -1123
rect 691 -1126 693 -1116
rect 695 -1126 705 -1116
rect 1053 -1120 1055 -1110
rect 1057 -1120 1067 -1110
rect 1147 -1113 1149 -1103
rect 1151 -1113 1161 -1103
rect -343 -1183 -341 -1173
rect -339 -1183 -329 -1173
rect -295 -1183 -294 -1173
rect -292 -1183 -290 -1173
rect -286 -1183 -284 -1173
rect -282 -1183 -281 -1173
rect -247 -1186 -245 -1176
rect -243 -1186 -233 -1176
rect 246 -1180 247 -1160
rect 249 -1180 257 -1160
rect 259 -1180 260 -1160
rect 295 -1177 297 -1167
rect 299 -1177 309 -1167
rect 751 -1169 752 -1149
rect 754 -1169 762 -1149
rect 764 -1169 765 -1149
rect 1207 -1156 1208 -1136
rect 1210 -1156 1218 -1136
rect 1220 -1156 1221 -1136
rect 1256 -1153 1258 -1143
rect 1260 -1153 1270 -1143
rect 800 -1166 802 -1156
rect 804 -1166 814 -1156
rect 92 -1200 94 -1190
rect 96 -1200 106 -1190
rect 140 -1200 141 -1190
rect 143 -1200 145 -1190
rect 149 -1200 151 -1190
rect 153 -1200 154 -1190
rect 188 -1203 190 -1193
rect 192 -1203 202 -1193
rect 597 -1189 599 -1179
rect 601 -1189 611 -1179
rect 645 -1189 646 -1179
rect 648 -1189 650 -1179
rect 654 -1189 656 -1179
rect 658 -1189 659 -1179
rect 693 -1192 695 -1182
rect 697 -1192 707 -1182
rect 1053 -1176 1055 -1166
rect 1057 -1176 1067 -1166
rect 1101 -1176 1102 -1166
rect 1104 -1176 1106 -1166
rect 1110 -1176 1112 -1166
rect 1114 -1176 1115 -1166
rect 1149 -1179 1151 -1169
rect 1153 -1179 1163 -1169
rect 1088 -1255 1089 -1245
rect 1091 -1255 1093 -1245
rect 1097 -1255 1099 -1245
rect 1101 -1255 1102 -1245
rect 637 -1279 638 -1269
rect 640 -1279 642 -1269
rect 646 -1279 648 -1269
rect 650 -1279 651 -1269
rect -327 -1292 -326 -1282
rect -324 -1292 -322 -1282
rect -318 -1292 -316 -1282
rect -314 -1292 -313 -1282
rect -279 -1295 -277 -1285
rect -275 -1295 -265 -1285
rect 143 -1291 144 -1281
rect 146 -1291 148 -1281
rect 152 -1291 154 -1281
rect 156 -1291 157 -1281
rect 191 -1294 193 -1284
rect 195 -1294 205 -1284
rect 685 -1282 687 -1272
rect 689 -1282 699 -1272
rect 1136 -1258 1138 -1248
rect 1140 -1258 1150 -1248
<< ndcontact >>
rect -347 -1147 -343 -1142
rect -329 -1147 -325 -1142
rect -301 -1146 -297 -1136
rect -283 -1146 -279 -1136
rect -253 -1140 -249 -1135
rect -235 -1140 -231 -1135
rect 1049 -1140 1053 -1135
rect 1067 -1140 1071 -1135
rect 1095 -1139 1099 -1129
rect 1113 -1139 1117 -1129
rect 1143 -1133 1147 -1128
rect 1161 -1133 1165 -1128
rect -347 -1203 -343 -1198
rect -329 -1203 -325 -1198
rect 88 -1164 92 -1159
rect 106 -1164 110 -1159
rect 134 -1163 138 -1153
rect 152 -1163 156 -1153
rect 182 -1157 186 -1152
rect 200 -1157 204 -1152
rect 593 -1153 597 -1148
rect 611 -1153 615 -1148
rect 639 -1152 643 -1142
rect 657 -1152 661 -1142
rect 687 -1146 691 -1141
rect 705 -1146 709 -1141
rect -144 -1180 -140 -1175
rect -126 -1180 -122 -1175
rect -193 -1188 -189 -1183
rect -185 -1188 -179 -1183
rect -175 -1188 -171 -1183
rect -299 -1212 -295 -1202
rect -281 -1212 -277 -1202
rect -251 -1206 -247 -1201
rect -233 -1206 -229 -1201
rect 88 -1220 92 -1215
rect 106 -1220 110 -1215
rect 291 -1197 295 -1192
rect 309 -1197 313 -1192
rect 242 -1205 246 -1200
rect 250 -1205 256 -1200
rect 260 -1205 264 -1200
rect 593 -1209 597 -1204
rect 611 -1209 615 -1204
rect 796 -1186 800 -1181
rect 814 -1186 818 -1181
rect 747 -1194 751 -1189
rect 755 -1194 761 -1189
rect 765 -1194 769 -1189
rect 1049 -1196 1053 -1191
rect 1067 -1196 1071 -1191
rect 1252 -1173 1256 -1168
rect 1270 -1173 1274 -1168
rect 1203 -1181 1207 -1176
rect 1211 -1181 1217 -1176
rect 1221 -1181 1225 -1176
rect 1097 -1205 1101 -1195
rect 1115 -1205 1119 -1195
rect 1145 -1199 1149 -1194
rect 1163 -1199 1167 -1194
rect 641 -1218 645 -1208
rect 659 -1218 663 -1208
rect 689 -1212 693 -1207
rect 707 -1212 711 -1207
rect 136 -1229 140 -1219
rect 154 -1229 158 -1219
rect 184 -1223 188 -1218
rect 202 -1223 206 -1218
rect 1084 -1284 1088 -1274
rect 1102 -1284 1106 -1274
rect 1132 -1278 1136 -1273
rect 1150 -1278 1154 -1273
rect 633 -1308 637 -1298
rect 651 -1308 655 -1298
rect 681 -1302 685 -1297
rect 699 -1302 703 -1297
rect -331 -1321 -327 -1311
rect -313 -1321 -309 -1311
rect -283 -1315 -279 -1310
rect -265 -1315 -261 -1310
rect 139 -1320 143 -1310
rect 157 -1320 161 -1310
rect 187 -1314 191 -1309
rect 205 -1314 209 -1309
<< pdcontact >>
rect -301 -1117 -297 -1107
rect -292 -1117 -288 -1107
rect -283 -1117 -279 -1107
rect 1095 -1110 1099 -1100
rect 1104 -1110 1108 -1100
rect 1113 -1110 1117 -1100
rect -347 -1127 -343 -1117
rect -329 -1127 -325 -1117
rect -253 -1120 -249 -1110
rect -235 -1120 -231 -1110
rect 639 -1123 643 -1113
rect 648 -1123 652 -1113
rect 657 -1123 661 -1113
rect 134 -1134 138 -1124
rect 143 -1134 147 -1124
rect 152 -1134 156 -1124
rect -193 -1163 -189 -1143
rect -175 -1163 -171 -1143
rect 88 -1144 92 -1134
rect 106 -1144 110 -1134
rect -144 -1160 -140 -1150
rect -126 -1160 -122 -1150
rect 182 -1137 186 -1127
rect 200 -1137 204 -1127
rect 593 -1133 597 -1123
rect 611 -1133 615 -1123
rect 687 -1126 691 -1116
rect 705 -1126 709 -1116
rect 1049 -1120 1053 -1110
rect 1067 -1120 1071 -1110
rect 1143 -1113 1147 -1103
rect 1161 -1113 1165 -1103
rect -347 -1183 -343 -1173
rect -329 -1183 -325 -1173
rect -299 -1183 -295 -1173
rect -290 -1183 -286 -1173
rect -281 -1183 -277 -1173
rect -251 -1186 -247 -1176
rect -233 -1186 -229 -1176
rect 242 -1180 246 -1160
rect 260 -1180 264 -1160
rect 291 -1177 295 -1167
rect 309 -1177 313 -1167
rect 747 -1169 751 -1149
rect 765 -1169 769 -1149
rect 1203 -1156 1207 -1136
rect 1221 -1156 1225 -1136
rect 1252 -1153 1256 -1143
rect 1270 -1153 1274 -1143
rect 796 -1166 800 -1156
rect 814 -1166 818 -1156
rect 88 -1200 92 -1190
rect 106 -1200 110 -1190
rect 136 -1200 140 -1190
rect 145 -1200 149 -1190
rect 154 -1200 158 -1190
rect 184 -1203 188 -1193
rect 202 -1203 206 -1193
rect 593 -1189 597 -1179
rect 611 -1189 615 -1179
rect 641 -1189 645 -1179
rect 650 -1189 654 -1179
rect 659 -1189 663 -1179
rect 689 -1192 693 -1182
rect 707 -1192 711 -1182
rect 1049 -1176 1053 -1166
rect 1067 -1176 1071 -1166
rect 1097 -1176 1101 -1166
rect 1106 -1176 1110 -1166
rect 1115 -1176 1119 -1166
rect 1145 -1179 1149 -1169
rect 1163 -1179 1167 -1169
rect 1084 -1255 1088 -1245
rect 1093 -1255 1097 -1245
rect 1102 -1255 1106 -1245
rect 633 -1279 637 -1269
rect 642 -1279 646 -1269
rect 651 -1279 655 -1269
rect -331 -1292 -327 -1282
rect -322 -1292 -318 -1282
rect -313 -1292 -309 -1282
rect -283 -1295 -279 -1285
rect -265 -1295 -261 -1285
rect 139 -1291 143 -1281
rect 148 -1291 152 -1281
rect 157 -1291 161 -1281
rect 187 -1294 191 -1284
rect 205 -1294 209 -1284
rect 681 -1282 685 -1272
rect 699 -1282 703 -1272
rect 1132 -1258 1136 -1248
rect 1150 -1258 1154 -1248
<< polysilicon >>
rect 1100 -1100 1102 -1097
rect 1110 -1100 1112 -1097
rect -296 -1107 -294 -1104
rect -286 -1107 -284 -1104
rect -341 -1117 -339 -1114
rect -247 -1110 -245 -1107
rect 1055 -1110 1057 -1107
rect 1149 -1103 1151 -1100
rect -341 -1142 -339 -1127
rect -296 -1136 -294 -1117
rect -286 -1136 -284 -1117
rect 644 -1113 646 -1110
rect 654 -1113 656 -1110
rect -247 -1135 -245 -1120
rect 139 -1124 141 -1121
rect 149 -1124 151 -1121
rect 599 -1123 601 -1120
rect 693 -1116 695 -1113
rect 94 -1134 96 -1131
rect 188 -1127 190 -1124
rect -247 -1143 -245 -1140
rect -188 -1143 -186 -1140
rect -178 -1143 -176 -1140
rect -341 -1150 -339 -1147
rect -296 -1149 -294 -1146
rect -286 -1149 -284 -1146
rect -138 -1150 -136 -1147
rect 94 -1159 96 -1144
rect 139 -1153 141 -1134
rect 149 -1153 151 -1134
rect 188 -1152 190 -1137
rect 599 -1148 601 -1133
rect 644 -1142 646 -1123
rect 654 -1142 656 -1123
rect 693 -1141 695 -1126
rect 1055 -1135 1057 -1120
rect 1100 -1129 1102 -1110
rect 1110 -1129 1112 -1110
rect 1149 -1128 1151 -1113
rect 1149 -1136 1151 -1133
rect 1208 -1136 1210 -1133
rect 1218 -1136 1220 -1133
rect -341 -1173 -339 -1170
rect -294 -1173 -292 -1170
rect -284 -1173 -282 -1170
rect -245 -1176 -243 -1173
rect -341 -1198 -339 -1183
rect -294 -1202 -292 -1183
rect -284 -1202 -282 -1183
rect -188 -1183 -186 -1163
rect -178 -1183 -176 -1163
rect -138 -1175 -136 -1160
rect 1055 -1143 1057 -1140
rect 1100 -1142 1102 -1139
rect 1110 -1142 1112 -1139
rect 693 -1149 695 -1146
rect 752 -1149 754 -1146
rect 762 -1149 764 -1146
rect 599 -1156 601 -1153
rect 644 -1155 646 -1152
rect 654 -1155 656 -1152
rect 188 -1160 190 -1157
rect 247 -1160 249 -1157
rect 257 -1160 259 -1157
rect 94 -1167 96 -1164
rect 139 -1166 141 -1163
rect 149 -1166 151 -1163
rect 297 -1167 299 -1164
rect 802 -1156 804 -1153
rect 1258 -1143 1260 -1140
rect 1055 -1166 1057 -1163
rect 1102 -1166 1104 -1163
rect 1112 -1166 1114 -1163
rect -138 -1183 -136 -1180
rect -245 -1201 -243 -1186
rect -188 -1191 -186 -1188
rect -178 -1191 -176 -1188
rect 94 -1190 96 -1187
rect 141 -1190 143 -1187
rect 151 -1190 153 -1187
rect 190 -1193 192 -1190
rect -341 -1206 -339 -1203
rect -245 -1209 -243 -1206
rect -294 -1215 -292 -1212
rect -284 -1215 -282 -1212
rect 94 -1215 96 -1200
rect 141 -1219 143 -1200
rect 151 -1219 153 -1200
rect 247 -1200 249 -1180
rect 257 -1200 259 -1180
rect 297 -1192 299 -1177
rect 599 -1179 601 -1176
rect 646 -1179 648 -1176
rect 656 -1179 658 -1176
rect 695 -1182 697 -1179
rect 297 -1200 299 -1197
rect 190 -1218 192 -1203
rect 599 -1204 601 -1189
rect 247 -1208 249 -1205
rect 257 -1208 259 -1205
rect 646 -1208 648 -1189
rect 656 -1208 658 -1189
rect 752 -1189 754 -1169
rect 762 -1189 764 -1169
rect 802 -1181 804 -1166
rect 1151 -1169 1153 -1166
rect 802 -1189 804 -1186
rect 695 -1207 697 -1192
rect 1055 -1191 1057 -1176
rect 752 -1197 754 -1194
rect 762 -1197 764 -1194
rect 1102 -1195 1104 -1176
rect 1112 -1195 1114 -1176
rect 1208 -1176 1210 -1156
rect 1218 -1176 1220 -1156
rect 1258 -1168 1260 -1153
rect 1258 -1176 1260 -1173
rect 1151 -1194 1153 -1179
rect 1208 -1184 1210 -1181
rect 1218 -1184 1220 -1181
rect 1055 -1199 1057 -1196
rect 1151 -1202 1153 -1199
rect 599 -1212 601 -1209
rect 1102 -1208 1104 -1205
rect 1112 -1208 1114 -1205
rect 695 -1215 697 -1212
rect 94 -1223 96 -1220
rect 646 -1221 648 -1218
rect 656 -1221 658 -1218
rect 190 -1226 192 -1223
rect 141 -1232 143 -1229
rect 151 -1232 153 -1229
rect 1089 -1245 1091 -1242
rect 1099 -1245 1101 -1242
rect 1138 -1248 1140 -1245
rect 638 -1269 640 -1266
rect 648 -1269 650 -1266
rect -326 -1282 -324 -1279
rect -316 -1282 -314 -1279
rect 144 -1281 146 -1278
rect 154 -1281 156 -1278
rect 687 -1272 689 -1269
rect -277 -1285 -275 -1282
rect -326 -1311 -324 -1292
rect -316 -1311 -314 -1292
rect 193 -1284 195 -1281
rect -277 -1310 -275 -1295
rect 144 -1310 146 -1291
rect 154 -1310 156 -1291
rect 193 -1309 195 -1294
rect 638 -1298 640 -1279
rect 648 -1298 650 -1279
rect 1089 -1274 1091 -1255
rect 1099 -1274 1101 -1255
rect 1138 -1273 1140 -1258
rect 687 -1297 689 -1282
rect 1138 -1281 1140 -1278
rect 1089 -1287 1091 -1284
rect 1099 -1287 1101 -1284
rect 687 -1305 689 -1302
rect -277 -1318 -275 -1315
rect 638 -1311 640 -1308
rect 648 -1311 650 -1308
rect 193 -1317 195 -1314
rect -326 -1324 -324 -1321
rect -316 -1324 -314 -1321
rect 144 -1323 146 -1320
rect 154 -1323 156 -1320
<< polycontact >>
rect -345 -1139 -341 -1135
rect -300 -1128 -296 -1124
rect -284 -1128 -280 -1124
rect -251 -1132 -247 -1128
rect 90 -1156 94 -1152
rect 135 -1145 139 -1141
rect 151 -1145 155 -1141
rect 184 -1149 188 -1145
rect 595 -1145 599 -1140
rect 640 -1134 644 -1130
rect 656 -1134 660 -1130
rect 689 -1138 693 -1134
rect 1051 -1132 1055 -1128
rect 1096 -1121 1100 -1117
rect 1112 -1121 1116 -1117
rect 1145 -1125 1149 -1121
rect -192 -1174 -188 -1170
rect -345 -1195 -341 -1191
rect -298 -1194 -294 -1190
rect -182 -1174 -178 -1170
rect -142 -1172 -138 -1168
rect -282 -1194 -278 -1190
rect -249 -1198 -245 -1194
rect 243 -1191 247 -1187
rect 90 -1212 94 -1208
rect 137 -1211 141 -1207
rect 253 -1191 257 -1187
rect 293 -1189 297 -1185
rect 748 -1180 752 -1176
rect 153 -1211 157 -1207
rect 186 -1215 190 -1211
rect 595 -1201 599 -1197
rect 642 -1200 646 -1196
rect 758 -1180 762 -1176
rect 798 -1178 802 -1174
rect 1204 -1167 1208 -1163
rect 1051 -1188 1055 -1184
rect 658 -1200 662 -1196
rect 691 -1204 695 -1200
rect 1098 -1187 1102 -1183
rect 1214 -1167 1218 -1163
rect 1254 -1165 1258 -1161
rect 1114 -1187 1118 -1183
rect 1147 -1191 1151 -1187
rect 1085 -1266 1089 -1262
rect -330 -1304 -326 -1299
rect -314 -1303 -310 -1299
rect -281 -1307 -277 -1303
rect 140 -1303 144 -1298
rect 634 -1291 638 -1286
rect 156 -1302 160 -1298
rect 189 -1306 193 -1302
rect 1101 -1266 1105 -1262
rect 1134 -1270 1138 -1266
rect 650 -1290 654 -1286
rect 683 -1294 687 -1290
<< metal1 >>
rect -307 -1102 -273 -1098
rect -301 -1107 -297 -1102
rect -283 -1107 -279 -1102
rect -259 -1104 -225 -1100
rect -353 -1111 -319 -1107
rect -347 -1117 -343 -1111
rect -253 -1110 -249 -1104
rect -377 -1135 -374 -1134
rect -329 -1135 -325 -1127
rect -316 -1128 -300 -1124
rect -316 -1135 -312 -1128
rect -292 -1131 -288 -1117
rect -280 -1128 -276 -1124
rect -235 -1128 -231 -1120
rect -292 -1132 -279 -1131
rect -266 -1132 -251 -1128
rect -235 -1132 -215 -1128
rect -292 -1135 -262 -1132
rect -235 -1135 -231 -1132
rect -377 -1139 -345 -1135
rect -329 -1139 -312 -1135
rect -283 -1136 -262 -1135
rect -329 -1142 -325 -1139
rect -253 -1146 -249 -1140
rect -347 -1153 -343 -1147
rect -301 -1150 -297 -1146
rect -259 -1149 -225 -1146
rect -307 -1153 -273 -1150
rect -353 -1156 -319 -1153
rect -353 -1167 -319 -1163
rect -347 -1173 -343 -1167
rect -305 -1168 -271 -1164
rect -299 -1173 -295 -1168
rect -281 -1173 -277 -1168
rect -257 -1170 -223 -1166
rect -220 -1170 -215 -1132
rect -199 -1135 -165 -1131
rect -193 -1143 -189 -1135
rect -150 -1144 -116 -1140
rect -144 -1150 -140 -1144
rect -251 -1176 -247 -1170
rect -220 -1174 -192 -1170
rect -175 -1176 -171 -1163
rect -126 -1168 -122 -1160
rect -111 -1168 -107 -1090
rect 1089 -1095 1123 -1091
rect 1095 -1100 1099 -1095
rect 1113 -1100 1117 -1095
rect 1137 -1097 1171 -1093
rect 1043 -1104 1077 -1100
rect 633 -1108 667 -1104
rect 639 -1113 643 -1108
rect 657 -1113 661 -1108
rect 681 -1110 715 -1106
rect 1049 -1110 1053 -1104
rect 1143 -1103 1147 -1097
rect 128 -1119 162 -1115
rect 587 -1117 621 -1113
rect 134 -1124 138 -1119
rect 152 -1124 156 -1119
rect 176 -1121 210 -1117
rect 82 -1128 116 -1124
rect 88 -1134 92 -1128
rect 182 -1127 186 -1121
rect 593 -1123 597 -1117
rect 687 -1116 691 -1110
rect 58 -1152 61 -1151
rect 106 -1152 110 -1144
rect 119 -1145 135 -1141
rect 119 -1152 123 -1145
rect 143 -1148 147 -1134
rect 155 -1145 159 -1141
rect 200 -1145 204 -1137
rect 563 -1145 595 -1140
rect 611 -1141 615 -1133
rect 624 -1134 640 -1130
rect 624 -1141 628 -1134
rect 648 -1137 652 -1123
rect 660 -1134 664 -1130
rect 705 -1134 709 -1126
rect 648 -1138 661 -1137
rect 674 -1138 689 -1134
rect 705 -1138 725 -1134
rect 648 -1141 678 -1138
rect 705 -1141 709 -1138
rect 611 -1145 628 -1141
rect 657 -1142 678 -1141
rect 143 -1149 156 -1148
rect 169 -1149 184 -1145
rect 200 -1149 220 -1145
rect 611 -1148 615 -1145
rect 143 -1152 173 -1149
rect 200 -1152 204 -1149
rect 58 -1156 90 -1152
rect 106 -1156 123 -1152
rect 152 -1153 173 -1152
rect 106 -1159 110 -1156
rect -162 -1172 -142 -1168
rect -126 -1172 -107 -1168
rect 182 -1163 186 -1157
rect 88 -1170 92 -1164
rect 134 -1167 138 -1163
rect 176 -1166 210 -1163
rect 128 -1170 162 -1167
rect -162 -1176 -158 -1172
rect -126 -1175 -122 -1172
rect -329 -1191 -325 -1183
rect -315 -1191 -298 -1190
rect -361 -1195 -345 -1191
rect -329 -1194 -298 -1191
rect -329 -1195 -314 -1194
rect -329 -1198 -325 -1195
rect -290 -1197 -286 -1183
rect -175 -1177 -158 -1176
rect -185 -1180 -158 -1177
rect -185 -1183 -179 -1180
rect -278 -1194 -274 -1190
rect -233 -1194 -229 -1186
rect -144 -1186 -140 -1180
rect -290 -1198 -277 -1197
rect -264 -1198 -249 -1194
rect -233 -1198 -219 -1194
rect -193 -1194 -189 -1188
rect -175 -1194 -171 -1188
rect -150 -1189 -116 -1186
rect -111 -1194 -107 -1172
rect 82 -1173 116 -1170
rect 82 -1184 116 -1180
rect 88 -1190 92 -1184
rect 130 -1185 164 -1181
rect 136 -1190 140 -1185
rect 154 -1190 158 -1185
rect 178 -1187 212 -1183
rect 215 -1187 220 -1149
rect 236 -1152 270 -1148
rect 242 -1160 246 -1152
rect 687 -1152 691 -1146
rect 285 -1161 319 -1157
rect 593 -1159 597 -1153
rect 639 -1156 643 -1152
rect 681 -1155 715 -1152
rect 633 -1159 667 -1156
rect 291 -1167 295 -1161
rect 587 -1162 621 -1159
rect -199 -1197 -165 -1194
rect -290 -1201 -260 -1198
rect -233 -1201 -229 -1198
rect 184 -1193 188 -1187
rect 215 -1191 243 -1187
rect 260 -1193 264 -1180
rect 309 -1185 313 -1177
rect 324 -1185 329 -1163
rect 587 -1173 621 -1169
rect 273 -1189 293 -1185
rect 309 -1189 329 -1185
rect 593 -1179 597 -1173
rect 635 -1174 669 -1170
rect 641 -1179 645 -1174
rect 659 -1179 663 -1174
rect 683 -1176 717 -1172
rect 720 -1176 725 -1138
rect 741 -1141 775 -1137
rect 747 -1149 751 -1141
rect 790 -1150 824 -1146
rect 796 -1156 800 -1150
rect 689 -1182 693 -1176
rect 720 -1180 748 -1176
rect 765 -1182 769 -1169
rect 814 -1174 818 -1166
rect 828 -1173 833 -1125
rect 1019 -1128 1022 -1127
rect 1067 -1128 1071 -1120
rect 1080 -1121 1096 -1117
rect 1080 -1128 1084 -1121
rect 1104 -1124 1108 -1110
rect 1116 -1121 1120 -1117
rect 1161 -1121 1165 -1113
rect 1104 -1125 1117 -1124
rect 1130 -1125 1145 -1121
rect 1161 -1125 1181 -1121
rect 1104 -1128 1134 -1125
rect 1161 -1128 1165 -1125
rect 1019 -1132 1051 -1128
rect 1067 -1132 1084 -1128
rect 1113 -1129 1134 -1128
rect 1067 -1135 1071 -1132
rect 1143 -1139 1147 -1133
rect 1049 -1146 1053 -1140
rect 1095 -1143 1099 -1139
rect 1137 -1142 1171 -1139
rect 1089 -1146 1123 -1143
rect 1043 -1149 1077 -1146
rect 1043 -1160 1077 -1156
rect 778 -1178 798 -1174
rect 814 -1178 828 -1174
rect 1049 -1166 1053 -1160
rect 1091 -1161 1125 -1157
rect 1097 -1166 1101 -1161
rect 1115 -1166 1119 -1161
rect 1139 -1163 1173 -1159
rect 1176 -1163 1181 -1125
rect 1197 -1128 1231 -1124
rect 1203 -1136 1207 -1128
rect 1246 -1137 1280 -1133
rect 1252 -1143 1256 -1137
rect 1145 -1169 1149 -1163
rect 1176 -1167 1204 -1163
rect 1221 -1169 1225 -1156
rect 1270 -1161 1274 -1153
rect 1285 -1161 1289 -1079
rect 1234 -1165 1254 -1161
rect 1270 -1165 1289 -1161
rect 1234 -1169 1238 -1165
rect 1270 -1168 1274 -1165
rect 778 -1182 782 -1178
rect 814 -1181 818 -1178
rect 273 -1193 277 -1189
rect 309 -1192 313 -1189
rect -281 -1202 -260 -1201
rect -347 -1209 -343 -1203
rect -353 -1212 -319 -1209
rect -251 -1212 -247 -1206
rect 106 -1208 110 -1200
rect 120 -1208 137 -1207
rect 74 -1212 90 -1208
rect 106 -1211 137 -1208
rect 106 -1212 121 -1211
rect -299 -1216 -295 -1212
rect -257 -1215 -223 -1212
rect 106 -1215 110 -1212
rect -305 -1219 -274 -1216
rect 145 -1214 149 -1200
rect 260 -1194 277 -1193
rect 250 -1197 277 -1194
rect 250 -1200 256 -1197
rect 157 -1211 161 -1207
rect 202 -1211 206 -1203
rect 291 -1203 295 -1197
rect 611 -1197 615 -1189
rect 625 -1197 642 -1196
rect 579 -1201 595 -1197
rect 611 -1200 642 -1197
rect 611 -1201 626 -1200
rect 145 -1215 158 -1214
rect 171 -1215 186 -1211
rect 202 -1215 216 -1211
rect 242 -1211 246 -1205
rect 260 -1211 264 -1205
rect 285 -1206 319 -1203
rect 611 -1204 615 -1201
rect 650 -1203 654 -1189
rect 765 -1183 782 -1182
rect 755 -1186 782 -1183
rect 755 -1189 761 -1186
rect 662 -1200 666 -1196
rect 707 -1200 711 -1192
rect 796 -1192 800 -1186
rect 1067 -1184 1071 -1176
rect 1081 -1184 1098 -1183
rect 1035 -1188 1051 -1184
rect 1067 -1187 1098 -1184
rect 1067 -1188 1082 -1187
rect 650 -1204 663 -1203
rect 676 -1204 691 -1200
rect 707 -1204 721 -1200
rect 747 -1200 751 -1194
rect 765 -1200 769 -1194
rect 790 -1195 824 -1192
rect 741 -1203 775 -1200
rect 650 -1207 680 -1204
rect 707 -1207 711 -1204
rect 659 -1208 680 -1207
rect 236 -1214 270 -1211
rect 593 -1215 597 -1209
rect 145 -1218 175 -1215
rect 202 -1218 206 -1215
rect 587 -1218 621 -1215
rect 689 -1218 693 -1212
rect 154 -1219 175 -1218
rect 88 -1226 92 -1220
rect 82 -1229 116 -1226
rect 641 -1222 645 -1218
rect 683 -1221 717 -1218
rect 184 -1229 188 -1223
rect 635 -1225 666 -1222
rect 136 -1233 140 -1229
rect 178 -1232 212 -1229
rect 130 -1236 161 -1233
rect 627 -1264 661 -1260
rect 1028 -1262 1035 -1188
rect 1067 -1191 1071 -1188
rect 1106 -1190 1110 -1176
rect 1221 -1170 1238 -1169
rect 1211 -1173 1238 -1170
rect 1211 -1176 1217 -1173
rect 1252 -1179 1256 -1173
rect 1118 -1187 1122 -1183
rect 1203 -1187 1207 -1181
rect 1221 -1187 1225 -1181
rect 1246 -1182 1280 -1179
rect 1106 -1191 1119 -1190
rect 1132 -1191 1147 -1187
rect 1197 -1190 1231 -1187
rect 1106 -1194 1136 -1191
rect 1115 -1195 1136 -1194
rect 1049 -1202 1053 -1196
rect 1043 -1205 1077 -1202
rect 1145 -1205 1149 -1199
rect 1097 -1209 1101 -1205
rect 1139 -1208 1173 -1205
rect 1091 -1212 1122 -1209
rect 1078 -1240 1112 -1236
rect 1084 -1245 1088 -1240
rect 1102 -1245 1106 -1240
rect 1126 -1242 1160 -1238
rect 1132 -1248 1136 -1242
rect 633 -1269 637 -1264
rect 651 -1269 655 -1264
rect 675 -1266 709 -1262
rect 1028 -1266 1085 -1262
rect -337 -1277 -303 -1273
rect -331 -1282 -327 -1277
rect -313 -1282 -309 -1277
rect -289 -1279 -255 -1275
rect 133 -1276 167 -1272
rect -283 -1285 -279 -1279
rect 139 -1281 143 -1276
rect 157 -1281 161 -1276
rect 181 -1278 215 -1274
rect -339 -1304 -330 -1299
rect -322 -1306 -318 -1292
rect 187 -1284 191 -1278
rect 681 -1272 685 -1266
rect 1093 -1269 1097 -1255
rect 1093 -1270 1106 -1269
rect 1115 -1270 1134 -1266
rect -265 -1303 -261 -1295
rect 98 -1303 140 -1298
rect -322 -1307 -309 -1306
rect -300 -1307 -281 -1303
rect -322 -1310 -297 -1307
rect -265 -1308 -251 -1303
rect 148 -1305 152 -1291
rect 603 -1291 634 -1286
rect 205 -1302 209 -1294
rect 642 -1293 646 -1279
rect 1093 -1273 1118 -1270
rect 1102 -1274 1118 -1273
rect 699 -1290 703 -1282
rect 1132 -1284 1136 -1278
rect 1084 -1288 1088 -1284
rect 1126 -1287 1160 -1284
rect 642 -1294 655 -1293
rect 664 -1294 683 -1290
rect 699 -1294 775 -1290
rect 1078 -1291 1112 -1288
rect 642 -1297 667 -1294
rect 699 -1297 703 -1294
rect 651 -1298 667 -1297
rect 148 -1306 161 -1305
rect 170 -1306 189 -1302
rect 205 -1306 229 -1302
rect -265 -1310 -261 -1308
rect 148 -1309 173 -1306
rect 205 -1309 209 -1306
rect 157 -1310 173 -1309
rect -313 -1311 -297 -1310
rect -283 -1321 -279 -1315
rect 681 -1308 685 -1302
rect 633 -1312 637 -1308
rect 675 -1311 709 -1308
rect 187 -1320 191 -1314
rect 627 -1315 661 -1312
rect -331 -1325 -327 -1321
rect -289 -1324 -255 -1321
rect 139 -1324 143 -1320
rect 181 -1323 215 -1320
rect -337 -1328 -303 -1325
rect 133 -1327 167 -1324
<< m2contact >>
rect -382 -1139 -377 -1134
rect -276 -1129 -271 -1124
rect 53 -1156 58 -1151
rect 159 -1146 164 -1141
rect 556 -1145 563 -1140
rect 664 -1135 669 -1130
rect -368 -1195 -361 -1190
rect -274 -1195 -269 -1190
rect -219 -1198 -214 -1193
rect 1014 -1132 1019 -1127
rect 1120 -1122 1125 -1117
rect 67 -1212 74 -1207
rect 161 -1212 166 -1207
rect 572 -1201 579 -1196
rect 216 -1215 221 -1210
rect 666 -1201 671 -1196
rect 1028 -1188 1035 -1183
rect 721 -1204 726 -1199
rect 1122 -1188 1127 -1183
rect -344 -1304 -339 -1299
rect 93 -1303 98 -1298
rect -251 -1308 -246 -1303
rect 598 -1291 603 -1286
<< metal2 >>
rect 1028 -1087 1129 -1084
rect -368 -1094 -267 -1091
rect -368 -1112 -361 -1094
rect -405 -1120 -361 -1112
rect -405 -1299 -397 -1120
rect -384 -1139 -382 -1134
rect -384 -1220 -377 -1139
rect -368 -1190 -361 -1120
rect -271 -1129 -267 -1094
rect 572 -1100 673 -1097
rect 67 -1111 168 -1108
rect 67 -1140 74 -1111
rect 27 -1146 74 -1140
rect 164 -1146 168 -1111
rect 572 -1129 579 -1100
rect 529 -1133 579 -1129
rect -184 -1174 -178 -1170
rect -219 -1177 -181 -1174
rect -274 -1220 -269 -1195
rect -219 -1193 -214 -1177
rect -384 -1226 -269 -1220
rect -301 -1299 -296 -1226
rect -405 -1304 -344 -1299
rect -310 -1303 -296 -1299
rect 27 -1298 33 -1146
rect 51 -1156 53 -1151
rect 51 -1237 58 -1156
rect 67 -1207 74 -1146
rect 251 -1191 257 -1187
rect 216 -1194 254 -1191
rect 161 -1237 166 -1212
rect 216 -1210 221 -1194
rect 51 -1243 166 -1237
rect 128 -1264 133 -1243
rect 128 -1268 175 -1264
rect 171 -1298 175 -1268
rect 529 -1286 533 -1133
rect 556 -1226 563 -1145
rect 572 -1196 579 -1133
rect 669 -1135 673 -1100
rect 1012 -1132 1014 -1127
rect 755 -1180 758 -1176
rect 721 -1183 758 -1180
rect 666 -1226 671 -1201
rect 721 -1199 726 -1183
rect 1012 -1213 1019 -1132
rect 1028 -1183 1035 -1087
rect 1125 -1122 1129 -1087
rect 1211 -1167 1214 -1163
rect 1177 -1170 1214 -1167
rect 1122 -1213 1127 -1188
rect 1163 -1187 1167 -1179
rect 1177 -1187 1182 -1170
rect 1163 -1191 1182 -1187
rect 1163 -1194 1167 -1191
rect 1012 -1219 1127 -1213
rect 556 -1232 671 -1226
rect 665 -1286 669 -1232
rect 1115 -1262 1119 -1219
rect 1105 -1266 1119 -1262
rect 1150 -1266 1154 -1258
rect 1150 -1270 1293 -1266
rect 1150 -1273 1154 -1270
rect 529 -1291 598 -1286
rect 654 -1290 669 -1286
rect 27 -1303 93 -1298
rect 160 -1302 175 -1298
rect -251 -1331 -246 -1308
<< m123contact >>
rect 828 -1178 833 -1173
<< metal3 >>
rect 833 -1178 847 -1173
rect 876 -1178 877 -1173
<< labels >>
rlabel polycontact -314 -1303 -310 -1299 1 b0
rlabel metal1 -259 -1308 -246 -1303 1 g0
rlabel ndcontact -265 -1315 -261 -1310 1 g0
rlabel pdcontact -265 -1295 -261 -1285 1 g0
rlabel ndiffusion -323 -1321 -317 -1311 1 and1nmg0
rlabel ndcontact -313 -1321 -309 -1311 1 g0n
rlabel pdcontact -322 -1292 -318 -1282 1 g0n
rlabel polycontact -281 -1307 -277 -1303 1 g0n
rlabel polycontact -330 -1304 -326 -1299 1 a0
rlabel ndcontact -283 -1315 -279 -1310 1 gnd
rlabel ndcontact -331 -1321 -327 -1311 1 gnd
rlabel metal1 -289 -1324 -255 -1321 1 gnd
rlabel metal1 -337 -1328 -303 -1325 1 gnd
rlabel metal1 -289 -1279 -255 -1275 1 vdd
rlabel metal1 -337 -1277 -303 -1273 1 vdd
rlabel pdcontact -283 -1295 -279 -1285 1 vdd
rlabel pdcontact -313 -1292 -309 -1282 1 vdd
rlabel pdcontact -331 -1292 -327 -1282 1 vdd
rlabel pdcontact -126 -1160 -122 -1150 1 p0
rlabel ndcontact -126 -1180 -122 -1175 1 p0
rlabel polycontact -142 -1172 -138 -1168 1 outnp0
rlabel ndcontact -185 -1188 -179 -1183 1 outnp0
rlabel pdcontact -175 -1163 -171 -1143 1 outnp0
rlabel pdiffusion -185 -1163 -179 -1143 1 orpmp0
rlabel polycontact -182 -1174 -178 -1170 1 or1p0
rlabel polycontact -192 -1174 -188 -1170 1 or2p0
rlabel ndcontact -235 -1140 -231 -1135 1 or2p0
rlabel pdcontact -235 -1120 -231 -1110 1 or2p0
rlabel pdcontact -233 -1186 -229 -1176 1 or1p0
rlabel ndcontact -233 -1206 -229 -1201 1 or1p0
rlabel polycontact -249 -1198 -245 -1194 1 and2np0
rlabel polycontact -251 -1132 -247 -1128 1 and1np0
rlabel pdcontact -292 -1117 -288 -1107 1 and1np0
rlabel ndiffusion -293 -1146 -287 -1136 1 and1nmp0
rlabel ndcontact -283 -1146 -279 -1136 1 and1np0
rlabel ndcontact -281 -1212 -277 -1202 1 and2np0
rlabel pdcontact -290 -1183 -286 -1173 1 and2np0
rlabel ndiffusion -291 -1212 -285 -1202 1 and2nmp0
rlabel metal1 -122 -1172 -111 -1168 1 p0
rlabel polycontact -282 -1194 -278 -1190 1 b0
rlabel polycontact -284 -1128 -280 -1124 1 a0
rlabel polycontact -300 -1128 -296 -1124 1 b0not
rlabel polycontact -298 -1194 -294 -1190 1 a0not
rlabel ndcontact -329 -1147 -325 -1142 1 b0not
rlabel ndcontact -329 -1203 -325 -1198 1 a0not
rlabel polycontact -345 -1195 -341 -1191 1 a0
rlabel polycontact -345 -1139 -341 -1135 1 b0
rlabel ndcontact -253 -1140 -249 -1135 1 gnd
rlabel metal1 -259 -1149 -225 -1146 1 gnd
rlabel metal1 -305 -1219 -274 -1216 1 gnd
rlabel pdcontact -329 -1183 -325 -1173 1 anot
rlabel pdcontact -329 -1127 -325 -1117 1 bnot
rlabel ndcontact -301 -1146 -297 -1136 1 gnd
rlabel ndcontact -347 -1147 -343 -1142 1 gnd
rlabel metal1 -307 -1153 -273 -1150 1 gnd
rlabel metal1 -353 -1156 -319 -1153 1 gnd
rlabel metal1 -353 -1212 -319 -1209 1 gnd
rlabel ndcontact -347 -1203 -343 -1198 1 gnd
rlabel ndcontact -251 -1206 -247 -1201 1 gnd
rlabel ndcontact -299 -1212 -295 -1202 1 gnd
rlabel metal1 -257 -1215 -223 -1212 1 gnd
rlabel metal1 -150 -1189 -116 -1186 1 gnd
rlabel ndcontact -144 -1180 -140 -1175 1 gnd
rlabel ndcontact -175 -1188 -171 -1183 1 gnd
rlabel ndcontact -193 -1188 -189 -1183 1 gnd
rlabel metal1 -199 -1197 -165 -1194 1 gnd
rlabel pdcontact -144 -1160 -140 -1150 1 vdd
rlabel metal1 -150 -1144 -116 -1140 1 vdd
rlabel pdcontact -193 -1163 -189 -1143 1 vdd
rlabel metal1 -199 -1135 -165 -1131 1 vdd
rlabel pdcontact -251 -1186 -247 -1176 1 vdd
rlabel metal1 -257 -1170 -223 -1166 1 vdd
rlabel pdcontact -281 -1183 -277 -1173 1 vdd
rlabel pdcontact -299 -1183 -295 -1173 1 vdd
rlabel metal1 -305 -1168 -271 -1164 1 vdd
rlabel pdcontact -347 -1183 -343 -1173 1 vdd
rlabel metal1 -353 -1167 -319 -1163 1 vdd
rlabel pdcontact -253 -1120 -249 -1110 1 vdd
rlabel metal1 -259 -1104 -225 -1100 5 vdd
rlabel pdcontact -283 -1117 -279 -1107 1 vdd
rlabel pdcontact -301 -1117 -297 -1107 1 vdd
rlabel metal1 -307 -1102 -273 -1098 5 vdd
rlabel pdcontact -347 -1127 -343 -1117 1 vdd
rlabel metal1 -353 -1111 -319 -1107 1 vdd
rlabel metal1 212 -1306 229 -1302 1 g1
rlabel ndcontact 205 -1314 209 -1309 1 g1
rlabel pdcontact 205 -1294 209 -1284 1 g1
rlabel polycontact 189 -1306 193 -1302 1 g1n
rlabel ndiffusion 147 -1320 153 -1310 1 and1nmg1
rlabel ndcontact 157 -1320 161 -1310 1 g1n
rlabel pdcontact 148 -1291 152 -1281 1 g1n
rlabel polycontact 156 -1302 160 -1298 1 b1
rlabel polycontact 140 -1303 144 -1298 1 a1
rlabel ndcontact 139 -1320 143 -1310 1 gnd
rlabel ndcontact 187 -1314 191 -1309 1 gnd
rlabel metal1 181 -1323 215 -1320 1 gnd
rlabel metal1 133 -1327 167 -1324 1 gnd
rlabel metal1 133 -1276 167 -1272 1 vdd
rlabel metal1 181 -1278 215 -1274 1 vdd
rlabel pdcontact 187 -1294 191 -1284 1 vdd
rlabel pdcontact 157 -1291 161 -1281 1 vdd
rlabel pdcontact 139 -1291 143 -1281 1 vdd
rlabel metal1 313 -1189 324 -1185 1 p1
rlabel ndcontact 309 -1197 313 -1192 1 p1
rlabel pdcontact 309 -1177 313 -1167 1 p1
rlabel polycontact 293 -1189 297 -1185 1 outnp1
rlabel ndcontact 250 -1205 256 -1200 1 outnp1
rlabel pdcontact 260 -1180 264 -1160 1 outnp1
rlabel pdiffusion 250 -1180 256 -1160 1 orpmp1
rlabel pdcontact 200 -1137 204 -1127 1 or2p1
rlabel ndcontact 200 -1157 204 -1152 1 or2p1
rlabel polycontact 243 -1191 247 -1187 1 or2p1
rlabel polycontact 253 -1191 257 -1187 1 or1p1
rlabel pdcontact 202 -1203 206 -1193 1 or1p1
rlabel ndcontact 202 -1223 206 -1218 1 or1p1
rlabel polycontact 186 -1215 190 -1211 1 and2np1
rlabel ndiffusion 144 -1229 150 -1219 1 and2nmp1
rlabel ndcontact 154 -1229 158 -1219 1 and2np1
rlabel pdcontact 145 -1200 149 -1190 1 and2np1
rlabel polycontact 153 -1211 157 -1207 1 b1
rlabel polycontact 151 -1145 155 -1141 1 a1
rlabel polycontact 184 -1149 188 -1145 1 and1np1
rlabel ndiffusion 142 -1163 148 -1153 1 and1nmp1
rlabel ndcontact 152 -1163 156 -1153 1 and1np1
rlabel pdcontact 143 -1134 147 -1124 1 and1np1
rlabel pdcontact 106 -1144 110 -1134 1 b1not
rlabel ndcontact 106 -1164 110 -1159 1 b1not
rlabel polycontact 135 -1145 139 -1141 1 b1not
rlabel polycontact 137 -1211 141 -1207 1 a1not
rlabel pdcontact 106 -1200 110 -1190 1 a1not
rlabel ndcontact 106 -1220 110 -1215 1 a1not
rlabel polycontact 90 -1212 94 -1208 1 a1
rlabel polycontact 90 -1156 94 -1152 1 b1
rlabel ndcontact 182 -1157 186 -1152 1 gnd
rlabel metal1 176 -1166 210 -1163 1 gnd
rlabel metal1 130 -1236 161 -1233 1 gnd
rlabel ndcontact 134 -1163 138 -1153 1 gnd
rlabel ndcontact 88 -1164 92 -1159 1 gnd
rlabel metal1 128 -1170 162 -1167 1 gnd
rlabel metal1 82 -1173 116 -1170 1 gnd
rlabel metal1 82 -1229 116 -1226 1 gnd
rlabel ndcontact 88 -1220 92 -1215 1 gnd
rlabel ndcontact 184 -1223 188 -1218 1 gnd
rlabel ndcontact 136 -1229 140 -1219 1 gnd
rlabel metal1 178 -1232 212 -1229 1 gnd
rlabel metal1 285 -1206 319 -1203 1 gnd
rlabel ndcontact 291 -1197 295 -1192 1 gnd
rlabel ndcontact 260 -1205 264 -1200 1 gnd
rlabel ndcontact 242 -1205 246 -1200 1 gnd
rlabel metal1 236 -1214 270 -1211 1 gnd
rlabel pdcontact 291 -1177 295 -1167 1 vdd
rlabel metal1 285 -1161 319 -1157 1 vdd
rlabel pdcontact 242 -1180 246 -1160 1 vdd
rlabel metal1 236 -1152 270 -1148 1 vdd
rlabel pdcontact 184 -1203 188 -1193 1 vdd
rlabel metal1 178 -1187 212 -1183 1 vdd
rlabel pdcontact 154 -1200 158 -1190 1 vdd
rlabel pdcontact 136 -1200 140 -1190 1 vdd
rlabel metal1 130 -1185 164 -1181 1 vdd
rlabel pdcontact 88 -1200 92 -1190 1 vdd
rlabel metal1 82 -1184 116 -1180 1 vdd
rlabel pdcontact 182 -1137 186 -1127 1 vdd
rlabel metal1 176 -1121 210 -1117 5 vdd
rlabel pdcontact 152 -1134 156 -1124 1 vdd
rlabel pdcontact 134 -1134 138 -1124 1 vdd
rlabel metal1 128 -1119 162 -1115 5 vdd
rlabel pdcontact 88 -1144 92 -1134 1 vdd
rlabel metal1 82 -1128 116 -1124 1 vdd
rlabel pdcontact 642 -1279 646 -1269 1 g2n
rlabel polycontact 758 -1180 762 -1176 1 or1p2
rlabel polycontact 650 -1290 654 -1286 1 b2
rlabel metal1 706 -1294 721 -1290 1 g2
rlabel pdcontact 699 -1282 703 -1272 1 g2
rlabel ndcontact 699 -1302 703 -1297 1 g2
rlabel ndiffusion 641 -1308 647 -1298 1 and1nmg2
rlabel polycontact 683 -1294 687 -1290 1 g2n
rlabel ndcontact 651 -1308 655 -1298 1 g2n
rlabel polycontact 634 -1291 638 -1286 1 a2
rlabel ndcontact 681 -1302 685 -1297 1 gnd
rlabel ndcontact 633 -1308 637 -1298 1 gnd
rlabel metal1 675 -1311 709 -1308 1 gnd
rlabel metal1 627 -1315 661 -1312 1 gnd
rlabel metal1 675 -1266 709 -1262 1 vdd
rlabel metal1 627 -1264 661 -1260 1 vdd
rlabel pdcontact 681 -1282 685 -1272 1 vdd
rlabel pdcontact 651 -1279 655 -1269 1 vdd
rlabel pdcontact 633 -1279 637 -1269 1 vdd
rlabel metal1 818 -1178 828 -1174 1 p2
rlabel pdcontact 814 -1166 818 -1156 1 p2
rlabel ndcontact 814 -1186 818 -1181 1 p2
rlabel polycontact 798 -1178 802 -1174 1 outnp2
rlabel pdcontact 765 -1169 769 -1149 1 outnp2
rlabel ndcontact 755 -1194 761 -1189 1 outnp2
rlabel pdiffusion 755 -1169 761 -1149 1 orpmp2
rlabel ndcontact 707 -1212 711 -1207 1 or1p2
rlabel pdcontact 707 -1192 711 -1182 1 or1p2
rlabel polycontact 748 -1180 752 -1176 1 or2p2
rlabel ndcontact 705 -1146 709 -1141 1 or2p2
rlabel pdcontact 705 -1126 709 -1116 1 or2p2
rlabel ndiffusion 647 -1152 653 -1142 1 and1nmp2
rlabel polycontact 656 -1134 660 -1130 1 a2
rlabel polycontact 689 -1138 693 -1134 1 and1np2
rlabel ndcontact 657 -1152 661 -1142 1 and1np2
rlabel pdcontact 648 -1123 652 -1113 1 and1np2
rlabel polycontact 640 -1134 644 -1130 1 b2not
rlabel pdcontact 611 -1133 615 -1123 1 b2not
rlabel ndcontact 611 -1153 615 -1148 1 b2not
rlabel polycontact 595 -1145 599 -1140 1 b2
rlabel ndiffusion 649 -1218 655 -1208 1 and2nmp2
rlabel polycontact 691 -1204 695 -1200 1 and2np2
rlabel ndcontact 659 -1218 663 -1208 1 and2np2
rlabel polycontact 658 -1200 662 -1196 1 b2
rlabel pdcontact 650 -1189 654 -1179 1 and2np2
rlabel polycontact 642 -1200 646 -1196 1 a2not
rlabel pdcontact 611 -1189 615 -1179 1 a2not
rlabel ndcontact 611 -1209 615 -1204 1 a2not
rlabel polycontact 595 -1201 599 -1197 1 a2
rlabel ndcontact 687 -1146 691 -1141 1 gnd
rlabel metal1 681 -1155 715 -1152 1 gnd
rlabel metal1 635 -1225 666 -1222 1 gnd
rlabel ndcontact 639 -1152 643 -1142 1 gnd
rlabel ndcontact 593 -1153 597 -1148 1 gnd
rlabel metal1 633 -1159 667 -1156 1 gnd
rlabel metal1 587 -1162 621 -1159 1 gnd
rlabel metal1 587 -1218 621 -1215 1 gnd
rlabel ndcontact 593 -1209 597 -1204 1 gnd
rlabel ndcontact 689 -1212 693 -1207 1 gnd
rlabel ndcontact 641 -1218 645 -1208 1 gnd
rlabel metal1 683 -1221 717 -1218 1 gnd
rlabel metal1 790 -1195 824 -1192 1 gnd
rlabel ndcontact 796 -1186 800 -1181 1 gnd
rlabel ndcontact 765 -1194 769 -1189 1 gnd
rlabel ndcontact 747 -1194 751 -1189 1 gnd
rlabel metal1 741 -1203 775 -1200 1 gnd
rlabel pdcontact 796 -1166 800 -1156 1 vdd
rlabel metal1 790 -1150 824 -1146 1 vdd
rlabel pdcontact 747 -1169 751 -1149 1 vdd
rlabel metal1 741 -1141 775 -1137 1 vdd
rlabel pdcontact 689 -1192 693 -1182 1 vdd
rlabel metal1 683 -1176 717 -1172 1 vdd
rlabel pdcontact 659 -1189 663 -1179 1 vdd
rlabel pdcontact 641 -1189 645 -1179 1 vdd
rlabel metal1 635 -1174 669 -1170 1 vdd
rlabel pdcontact 593 -1189 597 -1179 1 vdd
rlabel metal1 587 -1173 621 -1169 1 vdd
rlabel pdcontact 687 -1126 691 -1116 1 vdd
rlabel metal1 681 -1110 715 -1106 5 vdd
rlabel pdcontact 657 -1123 661 -1113 1 vdd
rlabel pdcontact 639 -1123 643 -1113 1 vdd
rlabel metal1 633 -1108 667 -1104 5 vdd
rlabel pdcontact 593 -1133 597 -1123 1 vdd
rlabel metal1 587 -1117 621 -1113 1 vdd
rlabel space 1214 -1170 1218 -1163 1 or1p3
rlabel ndcontact 1150 -1278 1154 -1273 1 g3
rlabel pdcontact 1150 -1258 1154 -1248 1 g3
rlabel metal2 1157 -1270 1174 -1266 1 g3
rlabel ndiffusion 1092 -1284 1098 -1274 1 and1nmg3
rlabel polycontact 1134 -1270 1138 -1266 1 g3n
rlabel ndcontact 1102 -1284 1106 -1274 1 g3n
rlabel pdcontact 1093 -1255 1097 -1245 1 g3n
rlabel polycontact 1085 -1266 1089 -1262 1 a3
rlabel ndcontact 1084 -1284 1088 -1274 1 gnd
rlabel ndcontact 1132 -1278 1136 -1273 1 gnd
rlabel metal1 1126 -1287 1160 -1284 1 gnd
rlabel metal1 1078 -1291 1112 -1288 1 gnd
rlabel metal1 1078 -1240 1112 -1236 1 vdd
rlabel metal1 1126 -1242 1160 -1238 1 vdd
rlabel pdcontact 1132 -1258 1136 -1248 1 vdd
rlabel pdcontact 1102 -1255 1106 -1245 1 vdd
rlabel pdcontact 1084 -1255 1088 -1245 1 vdd
rlabel metal1 1274 -1165 1285 -1161 1 p3
rlabel pdcontact 1270 -1153 1274 -1143 1 p3
rlabel ndcontact 1270 -1173 1274 -1168 1 p3
rlabel polycontact 1254 -1165 1258 -1161 1 outnp3
rlabel pdcontact 1221 -1156 1225 -1136 1 outnp3
rlabel ndcontact 1211 -1181 1217 -1176 1 outnp3
rlabel pdiffusion 1211 -1156 1217 -1136 1 orpmp3
rlabel ndcontact 1163 -1199 1167 -1194 1 or1p3
rlabel pdcontact 1163 -1179 1167 -1169 1 or1p3
rlabel ndcontact 1161 -1133 1165 -1128 1 or2p3
rlabel pdcontact 1161 -1113 1165 -1103 1 or2p3
rlabel polycontact 1114 -1187 1118 -1183 1 b3
rlabel ndiffusion 1105 -1205 1111 -1195 1 and2nmp3
rlabel polycontact 1147 -1191 1151 -1187 1 and2np3
rlabel ndcontact 1115 -1205 1119 -1195 1 and2np3
rlabel pdcontact 1106 -1176 1110 -1166 1 and2np3
rlabel ndiffusion 1103 -1139 1109 -1129 1 and1nmp3
rlabel polycontact 1112 -1121 1116 -1117 1 a3
rlabel polycontact 1145 -1125 1149 -1121 1 and1np3
rlabel ndcontact 1113 -1139 1117 -1129 1 and1np3
rlabel pdcontact 1104 -1110 1108 -1100 1 and1np3
rlabel polycontact 1098 -1187 1102 -1183 1 a3not
rlabel pdcontact 1067 -1176 1071 -1166 1 a3not
rlabel ndcontact 1067 -1196 1071 -1191 1 a3not
rlabel polycontact 1051 -1188 1055 -1184 1 a3
rlabel polycontact 1096 -1121 1100 -1117 1 b3not
rlabel pdcontact 1067 -1120 1071 -1110 1 b3not
rlabel ndcontact 1067 -1140 1071 -1135 1 b3not
rlabel polycontact 1051 -1132 1055 -1128 1 b3
rlabel ndcontact 1143 -1133 1147 -1128 1 gnd
rlabel metal1 1137 -1142 1171 -1139 1 gnd
rlabel metal1 1091 -1212 1122 -1209 1 gnd
rlabel ndcontact 1095 -1139 1099 -1129 1 gnd
rlabel ndcontact 1049 -1140 1053 -1135 1 gnd
rlabel metal1 1089 -1146 1123 -1143 1 gnd
rlabel metal1 1043 -1149 1077 -1146 1 gnd
rlabel metal1 1043 -1205 1077 -1202 1 gnd
rlabel ndcontact 1049 -1196 1053 -1191 1 gnd
rlabel ndcontact 1145 -1199 1149 -1194 1 gnd
rlabel ndcontact 1097 -1205 1101 -1195 1 gnd
rlabel metal1 1139 -1208 1173 -1205 1 gnd
rlabel metal1 1246 -1182 1280 -1179 1 gnd
rlabel ndcontact 1252 -1173 1256 -1168 1 gnd
rlabel ndcontact 1221 -1181 1225 -1176 1 gnd
rlabel ndcontact 1203 -1181 1207 -1176 1 gnd
rlabel metal1 1197 -1190 1231 -1187 1 gnd
rlabel pdcontact 1252 -1153 1256 -1143 1 vdd
rlabel metal1 1246 -1137 1280 -1133 1 vdd
rlabel pdcontact 1203 -1156 1207 -1136 1 vdd
rlabel metal1 1197 -1128 1231 -1124 1 vdd
rlabel pdcontact 1145 -1179 1149 -1169 1 vdd
rlabel metal1 1139 -1163 1173 -1159 1 vdd
rlabel pdcontact 1115 -1176 1119 -1166 1 vdd
rlabel pdcontact 1097 -1176 1101 -1166 1 vdd
rlabel metal1 1091 -1161 1125 -1157 1 vdd
rlabel pdcontact 1049 -1176 1053 -1166 1 vdd
rlabel metal1 1043 -1160 1077 -1156 1 vdd
rlabel pdcontact 1143 -1113 1147 -1103 1 vdd
rlabel metal1 1137 -1097 1171 -1093 5 vdd
rlabel pdcontact 1113 -1110 1117 -1100 1 vdd
rlabel pdcontact 1095 -1110 1099 -1100 1 vdd
rlabel metal1 1089 -1095 1123 -1091 5 vdd
rlabel pdcontact 1049 -1120 1053 -1110 1 vdd
rlabel metal1 1043 -1104 1077 -1100 1 vdd
rlabel metal1 1232 -1173 1238 -1169 1 outnp3
rlabel polycontact 1204 -1167 1208 -1163 1 or2p3
rlabel metal2 1177 -1170 1186 -1167 1 or1p3
rlabel metal1 1165 -1125 1174 -1121 1 or2p3
rlabel metal2 1171 -1191 1182 -1187 1 or1p3
rlabel polysilicon 1218 -1167 1220 -1163 1 or1p3
rlabel polycontact 1101 -1266 1105 -1262 1 b3
<< end >>
